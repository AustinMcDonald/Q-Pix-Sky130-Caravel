magic
tech sky130B
magscale 1 2
timestamp 1606595467
<< pwell >>
rect -5717 -1219 5717 1219
<< nmos >>
rect -5521 109 -5431 1009
rect -5373 109 -5283 1009
rect -5225 109 -5135 1009
rect -5077 109 -4987 1009
rect -4929 109 -4839 1009
rect -4781 109 -4691 1009
rect -4633 109 -4543 1009
rect -4485 109 -4395 1009
rect -4337 109 -4247 1009
rect -4189 109 -4099 1009
rect -4041 109 -3951 1009
rect -3893 109 -3803 1009
rect -3745 109 -3655 1009
rect -3597 109 -3507 1009
rect -3449 109 -3359 1009
rect -3301 109 -3211 1009
rect -3153 109 -3063 1009
rect -3005 109 -2915 1009
rect -2857 109 -2767 1009
rect -2709 109 -2619 1009
rect -2561 109 -2471 1009
rect -2413 109 -2323 1009
rect -2265 109 -2175 1009
rect -2117 109 -2027 1009
rect -1969 109 -1879 1009
rect -1821 109 -1731 1009
rect -1673 109 -1583 1009
rect -1525 109 -1435 1009
rect -1377 109 -1287 1009
rect -1229 109 -1139 1009
rect -1081 109 -991 1009
rect -933 109 -843 1009
rect -785 109 -695 1009
rect -637 109 -547 1009
rect -489 109 -399 1009
rect -341 109 -251 1009
rect -193 109 -103 1009
rect -45 109 45 1009
rect 103 109 193 1009
rect 251 109 341 1009
rect 399 109 489 1009
rect 547 109 637 1009
rect 695 109 785 1009
rect 843 109 933 1009
rect 991 109 1081 1009
rect 1139 109 1229 1009
rect 1287 109 1377 1009
rect 1435 109 1525 1009
rect 1583 109 1673 1009
rect 1731 109 1821 1009
rect 1879 109 1969 1009
rect 2027 109 2117 1009
rect 2175 109 2265 1009
rect 2323 109 2413 1009
rect 2471 109 2561 1009
rect 2619 109 2709 1009
rect 2767 109 2857 1009
rect 2915 109 3005 1009
rect 3063 109 3153 1009
rect 3211 109 3301 1009
rect 3359 109 3449 1009
rect 3507 109 3597 1009
rect 3655 109 3745 1009
rect 3803 109 3893 1009
rect 3951 109 4041 1009
rect 4099 109 4189 1009
rect 4247 109 4337 1009
rect 4395 109 4485 1009
rect 4543 109 4633 1009
rect 4691 109 4781 1009
rect 4839 109 4929 1009
rect 4987 109 5077 1009
rect 5135 109 5225 1009
rect 5283 109 5373 1009
rect 5431 109 5521 1009
rect -5521 -1009 -5431 -109
rect -5373 -1009 -5283 -109
rect -5225 -1009 -5135 -109
rect -5077 -1009 -4987 -109
rect -4929 -1009 -4839 -109
rect -4781 -1009 -4691 -109
rect -4633 -1009 -4543 -109
rect -4485 -1009 -4395 -109
rect -4337 -1009 -4247 -109
rect -4189 -1009 -4099 -109
rect -4041 -1009 -3951 -109
rect -3893 -1009 -3803 -109
rect -3745 -1009 -3655 -109
rect -3597 -1009 -3507 -109
rect -3449 -1009 -3359 -109
rect -3301 -1009 -3211 -109
rect -3153 -1009 -3063 -109
rect -3005 -1009 -2915 -109
rect -2857 -1009 -2767 -109
rect -2709 -1009 -2619 -109
rect -2561 -1009 -2471 -109
rect -2413 -1009 -2323 -109
rect -2265 -1009 -2175 -109
rect -2117 -1009 -2027 -109
rect -1969 -1009 -1879 -109
rect -1821 -1009 -1731 -109
rect -1673 -1009 -1583 -109
rect -1525 -1009 -1435 -109
rect -1377 -1009 -1287 -109
rect -1229 -1009 -1139 -109
rect -1081 -1009 -991 -109
rect -933 -1009 -843 -109
rect -785 -1009 -695 -109
rect -637 -1009 -547 -109
rect -489 -1009 -399 -109
rect -341 -1009 -251 -109
rect -193 -1009 -103 -109
rect -45 -1009 45 -109
rect 103 -1009 193 -109
rect 251 -1009 341 -109
rect 399 -1009 489 -109
rect 547 -1009 637 -109
rect 695 -1009 785 -109
rect 843 -1009 933 -109
rect 991 -1009 1081 -109
rect 1139 -1009 1229 -109
rect 1287 -1009 1377 -109
rect 1435 -1009 1525 -109
rect 1583 -1009 1673 -109
rect 1731 -1009 1821 -109
rect 1879 -1009 1969 -109
rect 2027 -1009 2117 -109
rect 2175 -1009 2265 -109
rect 2323 -1009 2413 -109
rect 2471 -1009 2561 -109
rect 2619 -1009 2709 -109
rect 2767 -1009 2857 -109
rect 2915 -1009 3005 -109
rect 3063 -1009 3153 -109
rect 3211 -1009 3301 -109
rect 3359 -1009 3449 -109
rect 3507 -1009 3597 -109
rect 3655 -1009 3745 -109
rect 3803 -1009 3893 -109
rect 3951 -1009 4041 -109
rect 4099 -1009 4189 -109
rect 4247 -1009 4337 -109
rect 4395 -1009 4485 -109
rect 4543 -1009 4633 -109
rect 4691 -1009 4781 -109
rect 4839 -1009 4929 -109
rect 4987 -1009 5077 -109
rect 5135 -1009 5225 -109
rect 5283 -1009 5373 -109
rect 5431 -1009 5521 -109
<< ndiff >>
rect -5579 997 -5521 1009
rect -5579 121 -5567 997
rect -5533 121 -5521 997
rect -5579 109 -5521 121
rect -5431 997 -5373 1009
rect -5431 121 -5419 997
rect -5385 121 -5373 997
rect -5431 109 -5373 121
rect -5283 997 -5225 1009
rect -5283 121 -5271 997
rect -5237 121 -5225 997
rect -5283 109 -5225 121
rect -5135 997 -5077 1009
rect -5135 121 -5123 997
rect -5089 121 -5077 997
rect -5135 109 -5077 121
rect -4987 997 -4929 1009
rect -4987 121 -4975 997
rect -4941 121 -4929 997
rect -4987 109 -4929 121
rect -4839 997 -4781 1009
rect -4839 121 -4827 997
rect -4793 121 -4781 997
rect -4839 109 -4781 121
rect -4691 997 -4633 1009
rect -4691 121 -4679 997
rect -4645 121 -4633 997
rect -4691 109 -4633 121
rect -4543 997 -4485 1009
rect -4543 121 -4531 997
rect -4497 121 -4485 997
rect -4543 109 -4485 121
rect -4395 997 -4337 1009
rect -4395 121 -4383 997
rect -4349 121 -4337 997
rect -4395 109 -4337 121
rect -4247 997 -4189 1009
rect -4247 121 -4235 997
rect -4201 121 -4189 997
rect -4247 109 -4189 121
rect -4099 997 -4041 1009
rect -4099 121 -4087 997
rect -4053 121 -4041 997
rect -4099 109 -4041 121
rect -3951 997 -3893 1009
rect -3951 121 -3939 997
rect -3905 121 -3893 997
rect -3951 109 -3893 121
rect -3803 997 -3745 1009
rect -3803 121 -3791 997
rect -3757 121 -3745 997
rect -3803 109 -3745 121
rect -3655 997 -3597 1009
rect -3655 121 -3643 997
rect -3609 121 -3597 997
rect -3655 109 -3597 121
rect -3507 997 -3449 1009
rect -3507 121 -3495 997
rect -3461 121 -3449 997
rect -3507 109 -3449 121
rect -3359 997 -3301 1009
rect -3359 121 -3347 997
rect -3313 121 -3301 997
rect -3359 109 -3301 121
rect -3211 997 -3153 1009
rect -3211 121 -3199 997
rect -3165 121 -3153 997
rect -3211 109 -3153 121
rect -3063 997 -3005 1009
rect -3063 121 -3051 997
rect -3017 121 -3005 997
rect -3063 109 -3005 121
rect -2915 997 -2857 1009
rect -2915 121 -2903 997
rect -2869 121 -2857 997
rect -2915 109 -2857 121
rect -2767 997 -2709 1009
rect -2767 121 -2755 997
rect -2721 121 -2709 997
rect -2767 109 -2709 121
rect -2619 997 -2561 1009
rect -2619 121 -2607 997
rect -2573 121 -2561 997
rect -2619 109 -2561 121
rect -2471 997 -2413 1009
rect -2471 121 -2459 997
rect -2425 121 -2413 997
rect -2471 109 -2413 121
rect -2323 997 -2265 1009
rect -2323 121 -2311 997
rect -2277 121 -2265 997
rect -2323 109 -2265 121
rect -2175 997 -2117 1009
rect -2175 121 -2163 997
rect -2129 121 -2117 997
rect -2175 109 -2117 121
rect -2027 997 -1969 1009
rect -2027 121 -2015 997
rect -1981 121 -1969 997
rect -2027 109 -1969 121
rect -1879 997 -1821 1009
rect -1879 121 -1867 997
rect -1833 121 -1821 997
rect -1879 109 -1821 121
rect -1731 997 -1673 1009
rect -1731 121 -1719 997
rect -1685 121 -1673 997
rect -1731 109 -1673 121
rect -1583 997 -1525 1009
rect -1583 121 -1571 997
rect -1537 121 -1525 997
rect -1583 109 -1525 121
rect -1435 997 -1377 1009
rect -1435 121 -1423 997
rect -1389 121 -1377 997
rect -1435 109 -1377 121
rect -1287 997 -1229 1009
rect -1287 121 -1275 997
rect -1241 121 -1229 997
rect -1287 109 -1229 121
rect -1139 997 -1081 1009
rect -1139 121 -1127 997
rect -1093 121 -1081 997
rect -1139 109 -1081 121
rect -991 997 -933 1009
rect -991 121 -979 997
rect -945 121 -933 997
rect -991 109 -933 121
rect -843 997 -785 1009
rect -843 121 -831 997
rect -797 121 -785 997
rect -843 109 -785 121
rect -695 997 -637 1009
rect -695 121 -683 997
rect -649 121 -637 997
rect -695 109 -637 121
rect -547 997 -489 1009
rect -547 121 -535 997
rect -501 121 -489 997
rect -547 109 -489 121
rect -399 997 -341 1009
rect -399 121 -387 997
rect -353 121 -341 997
rect -399 109 -341 121
rect -251 997 -193 1009
rect -251 121 -239 997
rect -205 121 -193 997
rect -251 109 -193 121
rect -103 997 -45 1009
rect -103 121 -91 997
rect -57 121 -45 997
rect -103 109 -45 121
rect 45 997 103 1009
rect 45 121 57 997
rect 91 121 103 997
rect 45 109 103 121
rect 193 997 251 1009
rect 193 121 205 997
rect 239 121 251 997
rect 193 109 251 121
rect 341 997 399 1009
rect 341 121 353 997
rect 387 121 399 997
rect 341 109 399 121
rect 489 997 547 1009
rect 489 121 501 997
rect 535 121 547 997
rect 489 109 547 121
rect 637 997 695 1009
rect 637 121 649 997
rect 683 121 695 997
rect 637 109 695 121
rect 785 997 843 1009
rect 785 121 797 997
rect 831 121 843 997
rect 785 109 843 121
rect 933 997 991 1009
rect 933 121 945 997
rect 979 121 991 997
rect 933 109 991 121
rect 1081 997 1139 1009
rect 1081 121 1093 997
rect 1127 121 1139 997
rect 1081 109 1139 121
rect 1229 997 1287 1009
rect 1229 121 1241 997
rect 1275 121 1287 997
rect 1229 109 1287 121
rect 1377 997 1435 1009
rect 1377 121 1389 997
rect 1423 121 1435 997
rect 1377 109 1435 121
rect 1525 997 1583 1009
rect 1525 121 1537 997
rect 1571 121 1583 997
rect 1525 109 1583 121
rect 1673 997 1731 1009
rect 1673 121 1685 997
rect 1719 121 1731 997
rect 1673 109 1731 121
rect 1821 997 1879 1009
rect 1821 121 1833 997
rect 1867 121 1879 997
rect 1821 109 1879 121
rect 1969 997 2027 1009
rect 1969 121 1981 997
rect 2015 121 2027 997
rect 1969 109 2027 121
rect 2117 997 2175 1009
rect 2117 121 2129 997
rect 2163 121 2175 997
rect 2117 109 2175 121
rect 2265 997 2323 1009
rect 2265 121 2277 997
rect 2311 121 2323 997
rect 2265 109 2323 121
rect 2413 997 2471 1009
rect 2413 121 2425 997
rect 2459 121 2471 997
rect 2413 109 2471 121
rect 2561 997 2619 1009
rect 2561 121 2573 997
rect 2607 121 2619 997
rect 2561 109 2619 121
rect 2709 997 2767 1009
rect 2709 121 2721 997
rect 2755 121 2767 997
rect 2709 109 2767 121
rect 2857 997 2915 1009
rect 2857 121 2869 997
rect 2903 121 2915 997
rect 2857 109 2915 121
rect 3005 997 3063 1009
rect 3005 121 3017 997
rect 3051 121 3063 997
rect 3005 109 3063 121
rect 3153 997 3211 1009
rect 3153 121 3165 997
rect 3199 121 3211 997
rect 3153 109 3211 121
rect 3301 997 3359 1009
rect 3301 121 3313 997
rect 3347 121 3359 997
rect 3301 109 3359 121
rect 3449 997 3507 1009
rect 3449 121 3461 997
rect 3495 121 3507 997
rect 3449 109 3507 121
rect 3597 997 3655 1009
rect 3597 121 3609 997
rect 3643 121 3655 997
rect 3597 109 3655 121
rect 3745 997 3803 1009
rect 3745 121 3757 997
rect 3791 121 3803 997
rect 3745 109 3803 121
rect 3893 997 3951 1009
rect 3893 121 3905 997
rect 3939 121 3951 997
rect 3893 109 3951 121
rect 4041 997 4099 1009
rect 4041 121 4053 997
rect 4087 121 4099 997
rect 4041 109 4099 121
rect 4189 997 4247 1009
rect 4189 121 4201 997
rect 4235 121 4247 997
rect 4189 109 4247 121
rect 4337 997 4395 1009
rect 4337 121 4349 997
rect 4383 121 4395 997
rect 4337 109 4395 121
rect 4485 997 4543 1009
rect 4485 121 4497 997
rect 4531 121 4543 997
rect 4485 109 4543 121
rect 4633 997 4691 1009
rect 4633 121 4645 997
rect 4679 121 4691 997
rect 4633 109 4691 121
rect 4781 997 4839 1009
rect 4781 121 4793 997
rect 4827 121 4839 997
rect 4781 109 4839 121
rect 4929 997 4987 1009
rect 4929 121 4941 997
rect 4975 121 4987 997
rect 4929 109 4987 121
rect 5077 997 5135 1009
rect 5077 121 5089 997
rect 5123 121 5135 997
rect 5077 109 5135 121
rect 5225 997 5283 1009
rect 5225 121 5237 997
rect 5271 121 5283 997
rect 5225 109 5283 121
rect 5373 997 5431 1009
rect 5373 121 5385 997
rect 5419 121 5431 997
rect 5373 109 5431 121
rect 5521 997 5579 1009
rect 5521 121 5533 997
rect 5567 121 5579 997
rect 5521 109 5579 121
rect -5579 -121 -5521 -109
rect -5579 -997 -5567 -121
rect -5533 -997 -5521 -121
rect -5579 -1009 -5521 -997
rect -5431 -121 -5373 -109
rect -5431 -997 -5419 -121
rect -5385 -997 -5373 -121
rect -5431 -1009 -5373 -997
rect -5283 -121 -5225 -109
rect -5283 -997 -5271 -121
rect -5237 -997 -5225 -121
rect -5283 -1009 -5225 -997
rect -5135 -121 -5077 -109
rect -5135 -997 -5123 -121
rect -5089 -997 -5077 -121
rect -5135 -1009 -5077 -997
rect -4987 -121 -4929 -109
rect -4987 -997 -4975 -121
rect -4941 -997 -4929 -121
rect -4987 -1009 -4929 -997
rect -4839 -121 -4781 -109
rect -4839 -997 -4827 -121
rect -4793 -997 -4781 -121
rect -4839 -1009 -4781 -997
rect -4691 -121 -4633 -109
rect -4691 -997 -4679 -121
rect -4645 -997 -4633 -121
rect -4691 -1009 -4633 -997
rect -4543 -121 -4485 -109
rect -4543 -997 -4531 -121
rect -4497 -997 -4485 -121
rect -4543 -1009 -4485 -997
rect -4395 -121 -4337 -109
rect -4395 -997 -4383 -121
rect -4349 -997 -4337 -121
rect -4395 -1009 -4337 -997
rect -4247 -121 -4189 -109
rect -4247 -997 -4235 -121
rect -4201 -997 -4189 -121
rect -4247 -1009 -4189 -997
rect -4099 -121 -4041 -109
rect -4099 -997 -4087 -121
rect -4053 -997 -4041 -121
rect -4099 -1009 -4041 -997
rect -3951 -121 -3893 -109
rect -3951 -997 -3939 -121
rect -3905 -997 -3893 -121
rect -3951 -1009 -3893 -997
rect -3803 -121 -3745 -109
rect -3803 -997 -3791 -121
rect -3757 -997 -3745 -121
rect -3803 -1009 -3745 -997
rect -3655 -121 -3597 -109
rect -3655 -997 -3643 -121
rect -3609 -997 -3597 -121
rect -3655 -1009 -3597 -997
rect -3507 -121 -3449 -109
rect -3507 -997 -3495 -121
rect -3461 -997 -3449 -121
rect -3507 -1009 -3449 -997
rect -3359 -121 -3301 -109
rect -3359 -997 -3347 -121
rect -3313 -997 -3301 -121
rect -3359 -1009 -3301 -997
rect -3211 -121 -3153 -109
rect -3211 -997 -3199 -121
rect -3165 -997 -3153 -121
rect -3211 -1009 -3153 -997
rect -3063 -121 -3005 -109
rect -3063 -997 -3051 -121
rect -3017 -997 -3005 -121
rect -3063 -1009 -3005 -997
rect -2915 -121 -2857 -109
rect -2915 -997 -2903 -121
rect -2869 -997 -2857 -121
rect -2915 -1009 -2857 -997
rect -2767 -121 -2709 -109
rect -2767 -997 -2755 -121
rect -2721 -997 -2709 -121
rect -2767 -1009 -2709 -997
rect -2619 -121 -2561 -109
rect -2619 -997 -2607 -121
rect -2573 -997 -2561 -121
rect -2619 -1009 -2561 -997
rect -2471 -121 -2413 -109
rect -2471 -997 -2459 -121
rect -2425 -997 -2413 -121
rect -2471 -1009 -2413 -997
rect -2323 -121 -2265 -109
rect -2323 -997 -2311 -121
rect -2277 -997 -2265 -121
rect -2323 -1009 -2265 -997
rect -2175 -121 -2117 -109
rect -2175 -997 -2163 -121
rect -2129 -997 -2117 -121
rect -2175 -1009 -2117 -997
rect -2027 -121 -1969 -109
rect -2027 -997 -2015 -121
rect -1981 -997 -1969 -121
rect -2027 -1009 -1969 -997
rect -1879 -121 -1821 -109
rect -1879 -997 -1867 -121
rect -1833 -997 -1821 -121
rect -1879 -1009 -1821 -997
rect -1731 -121 -1673 -109
rect -1731 -997 -1719 -121
rect -1685 -997 -1673 -121
rect -1731 -1009 -1673 -997
rect -1583 -121 -1525 -109
rect -1583 -997 -1571 -121
rect -1537 -997 -1525 -121
rect -1583 -1009 -1525 -997
rect -1435 -121 -1377 -109
rect -1435 -997 -1423 -121
rect -1389 -997 -1377 -121
rect -1435 -1009 -1377 -997
rect -1287 -121 -1229 -109
rect -1287 -997 -1275 -121
rect -1241 -997 -1229 -121
rect -1287 -1009 -1229 -997
rect -1139 -121 -1081 -109
rect -1139 -997 -1127 -121
rect -1093 -997 -1081 -121
rect -1139 -1009 -1081 -997
rect -991 -121 -933 -109
rect -991 -997 -979 -121
rect -945 -997 -933 -121
rect -991 -1009 -933 -997
rect -843 -121 -785 -109
rect -843 -997 -831 -121
rect -797 -997 -785 -121
rect -843 -1009 -785 -997
rect -695 -121 -637 -109
rect -695 -997 -683 -121
rect -649 -997 -637 -121
rect -695 -1009 -637 -997
rect -547 -121 -489 -109
rect -547 -997 -535 -121
rect -501 -997 -489 -121
rect -547 -1009 -489 -997
rect -399 -121 -341 -109
rect -399 -997 -387 -121
rect -353 -997 -341 -121
rect -399 -1009 -341 -997
rect -251 -121 -193 -109
rect -251 -997 -239 -121
rect -205 -997 -193 -121
rect -251 -1009 -193 -997
rect -103 -121 -45 -109
rect -103 -997 -91 -121
rect -57 -997 -45 -121
rect -103 -1009 -45 -997
rect 45 -121 103 -109
rect 45 -997 57 -121
rect 91 -997 103 -121
rect 45 -1009 103 -997
rect 193 -121 251 -109
rect 193 -997 205 -121
rect 239 -997 251 -121
rect 193 -1009 251 -997
rect 341 -121 399 -109
rect 341 -997 353 -121
rect 387 -997 399 -121
rect 341 -1009 399 -997
rect 489 -121 547 -109
rect 489 -997 501 -121
rect 535 -997 547 -121
rect 489 -1009 547 -997
rect 637 -121 695 -109
rect 637 -997 649 -121
rect 683 -997 695 -121
rect 637 -1009 695 -997
rect 785 -121 843 -109
rect 785 -997 797 -121
rect 831 -997 843 -121
rect 785 -1009 843 -997
rect 933 -121 991 -109
rect 933 -997 945 -121
rect 979 -997 991 -121
rect 933 -1009 991 -997
rect 1081 -121 1139 -109
rect 1081 -997 1093 -121
rect 1127 -997 1139 -121
rect 1081 -1009 1139 -997
rect 1229 -121 1287 -109
rect 1229 -997 1241 -121
rect 1275 -997 1287 -121
rect 1229 -1009 1287 -997
rect 1377 -121 1435 -109
rect 1377 -997 1389 -121
rect 1423 -997 1435 -121
rect 1377 -1009 1435 -997
rect 1525 -121 1583 -109
rect 1525 -997 1537 -121
rect 1571 -997 1583 -121
rect 1525 -1009 1583 -997
rect 1673 -121 1731 -109
rect 1673 -997 1685 -121
rect 1719 -997 1731 -121
rect 1673 -1009 1731 -997
rect 1821 -121 1879 -109
rect 1821 -997 1833 -121
rect 1867 -997 1879 -121
rect 1821 -1009 1879 -997
rect 1969 -121 2027 -109
rect 1969 -997 1981 -121
rect 2015 -997 2027 -121
rect 1969 -1009 2027 -997
rect 2117 -121 2175 -109
rect 2117 -997 2129 -121
rect 2163 -997 2175 -121
rect 2117 -1009 2175 -997
rect 2265 -121 2323 -109
rect 2265 -997 2277 -121
rect 2311 -997 2323 -121
rect 2265 -1009 2323 -997
rect 2413 -121 2471 -109
rect 2413 -997 2425 -121
rect 2459 -997 2471 -121
rect 2413 -1009 2471 -997
rect 2561 -121 2619 -109
rect 2561 -997 2573 -121
rect 2607 -997 2619 -121
rect 2561 -1009 2619 -997
rect 2709 -121 2767 -109
rect 2709 -997 2721 -121
rect 2755 -997 2767 -121
rect 2709 -1009 2767 -997
rect 2857 -121 2915 -109
rect 2857 -997 2869 -121
rect 2903 -997 2915 -121
rect 2857 -1009 2915 -997
rect 3005 -121 3063 -109
rect 3005 -997 3017 -121
rect 3051 -997 3063 -121
rect 3005 -1009 3063 -997
rect 3153 -121 3211 -109
rect 3153 -997 3165 -121
rect 3199 -997 3211 -121
rect 3153 -1009 3211 -997
rect 3301 -121 3359 -109
rect 3301 -997 3313 -121
rect 3347 -997 3359 -121
rect 3301 -1009 3359 -997
rect 3449 -121 3507 -109
rect 3449 -997 3461 -121
rect 3495 -997 3507 -121
rect 3449 -1009 3507 -997
rect 3597 -121 3655 -109
rect 3597 -997 3609 -121
rect 3643 -997 3655 -121
rect 3597 -1009 3655 -997
rect 3745 -121 3803 -109
rect 3745 -997 3757 -121
rect 3791 -997 3803 -121
rect 3745 -1009 3803 -997
rect 3893 -121 3951 -109
rect 3893 -997 3905 -121
rect 3939 -997 3951 -121
rect 3893 -1009 3951 -997
rect 4041 -121 4099 -109
rect 4041 -997 4053 -121
rect 4087 -997 4099 -121
rect 4041 -1009 4099 -997
rect 4189 -121 4247 -109
rect 4189 -997 4201 -121
rect 4235 -997 4247 -121
rect 4189 -1009 4247 -997
rect 4337 -121 4395 -109
rect 4337 -997 4349 -121
rect 4383 -997 4395 -121
rect 4337 -1009 4395 -997
rect 4485 -121 4543 -109
rect 4485 -997 4497 -121
rect 4531 -997 4543 -121
rect 4485 -1009 4543 -997
rect 4633 -121 4691 -109
rect 4633 -997 4645 -121
rect 4679 -997 4691 -121
rect 4633 -1009 4691 -997
rect 4781 -121 4839 -109
rect 4781 -997 4793 -121
rect 4827 -997 4839 -121
rect 4781 -1009 4839 -997
rect 4929 -121 4987 -109
rect 4929 -997 4941 -121
rect 4975 -997 4987 -121
rect 4929 -1009 4987 -997
rect 5077 -121 5135 -109
rect 5077 -997 5089 -121
rect 5123 -997 5135 -121
rect 5077 -1009 5135 -997
rect 5225 -121 5283 -109
rect 5225 -997 5237 -121
rect 5271 -997 5283 -121
rect 5225 -1009 5283 -997
rect 5373 -121 5431 -109
rect 5373 -997 5385 -121
rect 5419 -997 5431 -121
rect 5373 -1009 5431 -997
rect 5521 -121 5579 -109
rect 5521 -997 5533 -121
rect 5567 -997 5579 -121
rect 5521 -1009 5579 -997
<< ndiffc >>
rect -5567 121 -5533 997
rect -5419 121 -5385 997
rect -5271 121 -5237 997
rect -5123 121 -5089 997
rect -4975 121 -4941 997
rect -4827 121 -4793 997
rect -4679 121 -4645 997
rect -4531 121 -4497 997
rect -4383 121 -4349 997
rect -4235 121 -4201 997
rect -4087 121 -4053 997
rect -3939 121 -3905 997
rect -3791 121 -3757 997
rect -3643 121 -3609 997
rect -3495 121 -3461 997
rect -3347 121 -3313 997
rect -3199 121 -3165 997
rect -3051 121 -3017 997
rect -2903 121 -2869 997
rect -2755 121 -2721 997
rect -2607 121 -2573 997
rect -2459 121 -2425 997
rect -2311 121 -2277 997
rect -2163 121 -2129 997
rect -2015 121 -1981 997
rect -1867 121 -1833 997
rect -1719 121 -1685 997
rect -1571 121 -1537 997
rect -1423 121 -1389 997
rect -1275 121 -1241 997
rect -1127 121 -1093 997
rect -979 121 -945 997
rect -831 121 -797 997
rect -683 121 -649 997
rect -535 121 -501 997
rect -387 121 -353 997
rect -239 121 -205 997
rect -91 121 -57 997
rect 57 121 91 997
rect 205 121 239 997
rect 353 121 387 997
rect 501 121 535 997
rect 649 121 683 997
rect 797 121 831 997
rect 945 121 979 997
rect 1093 121 1127 997
rect 1241 121 1275 997
rect 1389 121 1423 997
rect 1537 121 1571 997
rect 1685 121 1719 997
rect 1833 121 1867 997
rect 1981 121 2015 997
rect 2129 121 2163 997
rect 2277 121 2311 997
rect 2425 121 2459 997
rect 2573 121 2607 997
rect 2721 121 2755 997
rect 2869 121 2903 997
rect 3017 121 3051 997
rect 3165 121 3199 997
rect 3313 121 3347 997
rect 3461 121 3495 997
rect 3609 121 3643 997
rect 3757 121 3791 997
rect 3905 121 3939 997
rect 4053 121 4087 997
rect 4201 121 4235 997
rect 4349 121 4383 997
rect 4497 121 4531 997
rect 4645 121 4679 997
rect 4793 121 4827 997
rect 4941 121 4975 997
rect 5089 121 5123 997
rect 5237 121 5271 997
rect 5385 121 5419 997
rect 5533 121 5567 997
rect -5567 -997 -5533 -121
rect -5419 -997 -5385 -121
rect -5271 -997 -5237 -121
rect -5123 -997 -5089 -121
rect -4975 -997 -4941 -121
rect -4827 -997 -4793 -121
rect -4679 -997 -4645 -121
rect -4531 -997 -4497 -121
rect -4383 -997 -4349 -121
rect -4235 -997 -4201 -121
rect -4087 -997 -4053 -121
rect -3939 -997 -3905 -121
rect -3791 -997 -3757 -121
rect -3643 -997 -3609 -121
rect -3495 -997 -3461 -121
rect -3347 -997 -3313 -121
rect -3199 -997 -3165 -121
rect -3051 -997 -3017 -121
rect -2903 -997 -2869 -121
rect -2755 -997 -2721 -121
rect -2607 -997 -2573 -121
rect -2459 -997 -2425 -121
rect -2311 -997 -2277 -121
rect -2163 -997 -2129 -121
rect -2015 -997 -1981 -121
rect -1867 -997 -1833 -121
rect -1719 -997 -1685 -121
rect -1571 -997 -1537 -121
rect -1423 -997 -1389 -121
rect -1275 -997 -1241 -121
rect -1127 -997 -1093 -121
rect -979 -997 -945 -121
rect -831 -997 -797 -121
rect -683 -997 -649 -121
rect -535 -997 -501 -121
rect -387 -997 -353 -121
rect -239 -997 -205 -121
rect -91 -997 -57 -121
rect 57 -997 91 -121
rect 205 -997 239 -121
rect 353 -997 387 -121
rect 501 -997 535 -121
rect 649 -997 683 -121
rect 797 -997 831 -121
rect 945 -997 979 -121
rect 1093 -997 1127 -121
rect 1241 -997 1275 -121
rect 1389 -997 1423 -121
rect 1537 -997 1571 -121
rect 1685 -997 1719 -121
rect 1833 -997 1867 -121
rect 1981 -997 2015 -121
rect 2129 -997 2163 -121
rect 2277 -997 2311 -121
rect 2425 -997 2459 -121
rect 2573 -997 2607 -121
rect 2721 -997 2755 -121
rect 2869 -997 2903 -121
rect 3017 -997 3051 -121
rect 3165 -997 3199 -121
rect 3313 -997 3347 -121
rect 3461 -997 3495 -121
rect 3609 -997 3643 -121
rect 3757 -997 3791 -121
rect 3905 -997 3939 -121
rect 4053 -997 4087 -121
rect 4201 -997 4235 -121
rect 4349 -997 4383 -121
rect 4497 -997 4531 -121
rect 4645 -997 4679 -121
rect 4793 -997 4827 -121
rect 4941 -997 4975 -121
rect 5089 -997 5123 -121
rect 5237 -997 5271 -121
rect 5385 -997 5419 -121
rect 5533 -997 5567 -121
<< psubdiff >>
rect -5681 1149 -5585 1183
rect 5585 1149 5681 1183
rect -5681 1087 -5647 1149
rect 5647 1087 5681 1149
rect -5681 -1149 -5647 -1087
rect 5647 -1149 5681 -1087
rect -5681 -1183 -5585 -1149
rect 5585 -1183 5681 -1149
<< psubdiffcont >>
rect -5585 1149 5585 1183
rect -5681 -1087 -5647 1087
rect 5647 -1087 5681 1087
rect -5585 -1183 5585 -1149
<< poly >>
rect -5521 1081 -5431 1097
rect -5521 1047 -5505 1081
rect -5447 1047 -5431 1081
rect -5521 1009 -5431 1047
rect -5373 1081 -5283 1097
rect -5373 1047 -5357 1081
rect -5299 1047 -5283 1081
rect -5373 1009 -5283 1047
rect -5225 1081 -5135 1097
rect -5225 1047 -5209 1081
rect -5151 1047 -5135 1081
rect -5225 1009 -5135 1047
rect -5077 1081 -4987 1097
rect -5077 1047 -5061 1081
rect -5003 1047 -4987 1081
rect -5077 1009 -4987 1047
rect -4929 1081 -4839 1097
rect -4929 1047 -4913 1081
rect -4855 1047 -4839 1081
rect -4929 1009 -4839 1047
rect -4781 1081 -4691 1097
rect -4781 1047 -4765 1081
rect -4707 1047 -4691 1081
rect -4781 1009 -4691 1047
rect -4633 1081 -4543 1097
rect -4633 1047 -4617 1081
rect -4559 1047 -4543 1081
rect -4633 1009 -4543 1047
rect -4485 1081 -4395 1097
rect -4485 1047 -4469 1081
rect -4411 1047 -4395 1081
rect -4485 1009 -4395 1047
rect -4337 1081 -4247 1097
rect -4337 1047 -4321 1081
rect -4263 1047 -4247 1081
rect -4337 1009 -4247 1047
rect -4189 1081 -4099 1097
rect -4189 1047 -4173 1081
rect -4115 1047 -4099 1081
rect -4189 1009 -4099 1047
rect -4041 1081 -3951 1097
rect -4041 1047 -4025 1081
rect -3967 1047 -3951 1081
rect -4041 1009 -3951 1047
rect -3893 1081 -3803 1097
rect -3893 1047 -3877 1081
rect -3819 1047 -3803 1081
rect -3893 1009 -3803 1047
rect -3745 1081 -3655 1097
rect -3745 1047 -3729 1081
rect -3671 1047 -3655 1081
rect -3745 1009 -3655 1047
rect -3597 1081 -3507 1097
rect -3597 1047 -3581 1081
rect -3523 1047 -3507 1081
rect -3597 1009 -3507 1047
rect -3449 1081 -3359 1097
rect -3449 1047 -3433 1081
rect -3375 1047 -3359 1081
rect -3449 1009 -3359 1047
rect -3301 1081 -3211 1097
rect -3301 1047 -3285 1081
rect -3227 1047 -3211 1081
rect -3301 1009 -3211 1047
rect -3153 1081 -3063 1097
rect -3153 1047 -3137 1081
rect -3079 1047 -3063 1081
rect -3153 1009 -3063 1047
rect -3005 1081 -2915 1097
rect -3005 1047 -2989 1081
rect -2931 1047 -2915 1081
rect -3005 1009 -2915 1047
rect -2857 1081 -2767 1097
rect -2857 1047 -2841 1081
rect -2783 1047 -2767 1081
rect -2857 1009 -2767 1047
rect -2709 1081 -2619 1097
rect -2709 1047 -2693 1081
rect -2635 1047 -2619 1081
rect -2709 1009 -2619 1047
rect -2561 1081 -2471 1097
rect -2561 1047 -2545 1081
rect -2487 1047 -2471 1081
rect -2561 1009 -2471 1047
rect -2413 1081 -2323 1097
rect -2413 1047 -2397 1081
rect -2339 1047 -2323 1081
rect -2413 1009 -2323 1047
rect -2265 1081 -2175 1097
rect -2265 1047 -2249 1081
rect -2191 1047 -2175 1081
rect -2265 1009 -2175 1047
rect -2117 1081 -2027 1097
rect -2117 1047 -2101 1081
rect -2043 1047 -2027 1081
rect -2117 1009 -2027 1047
rect -1969 1081 -1879 1097
rect -1969 1047 -1953 1081
rect -1895 1047 -1879 1081
rect -1969 1009 -1879 1047
rect -1821 1081 -1731 1097
rect -1821 1047 -1805 1081
rect -1747 1047 -1731 1081
rect -1821 1009 -1731 1047
rect -1673 1081 -1583 1097
rect -1673 1047 -1657 1081
rect -1599 1047 -1583 1081
rect -1673 1009 -1583 1047
rect -1525 1081 -1435 1097
rect -1525 1047 -1509 1081
rect -1451 1047 -1435 1081
rect -1525 1009 -1435 1047
rect -1377 1081 -1287 1097
rect -1377 1047 -1361 1081
rect -1303 1047 -1287 1081
rect -1377 1009 -1287 1047
rect -1229 1081 -1139 1097
rect -1229 1047 -1213 1081
rect -1155 1047 -1139 1081
rect -1229 1009 -1139 1047
rect -1081 1081 -991 1097
rect -1081 1047 -1065 1081
rect -1007 1047 -991 1081
rect -1081 1009 -991 1047
rect -933 1081 -843 1097
rect -933 1047 -917 1081
rect -859 1047 -843 1081
rect -933 1009 -843 1047
rect -785 1081 -695 1097
rect -785 1047 -769 1081
rect -711 1047 -695 1081
rect -785 1009 -695 1047
rect -637 1081 -547 1097
rect -637 1047 -621 1081
rect -563 1047 -547 1081
rect -637 1009 -547 1047
rect -489 1081 -399 1097
rect -489 1047 -473 1081
rect -415 1047 -399 1081
rect -489 1009 -399 1047
rect -341 1081 -251 1097
rect -341 1047 -325 1081
rect -267 1047 -251 1081
rect -341 1009 -251 1047
rect -193 1081 -103 1097
rect -193 1047 -177 1081
rect -119 1047 -103 1081
rect -193 1009 -103 1047
rect -45 1081 45 1097
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect -45 1009 45 1047
rect 103 1081 193 1097
rect 103 1047 119 1081
rect 177 1047 193 1081
rect 103 1009 193 1047
rect 251 1081 341 1097
rect 251 1047 267 1081
rect 325 1047 341 1081
rect 251 1009 341 1047
rect 399 1081 489 1097
rect 399 1047 415 1081
rect 473 1047 489 1081
rect 399 1009 489 1047
rect 547 1081 637 1097
rect 547 1047 563 1081
rect 621 1047 637 1081
rect 547 1009 637 1047
rect 695 1081 785 1097
rect 695 1047 711 1081
rect 769 1047 785 1081
rect 695 1009 785 1047
rect 843 1081 933 1097
rect 843 1047 859 1081
rect 917 1047 933 1081
rect 843 1009 933 1047
rect 991 1081 1081 1097
rect 991 1047 1007 1081
rect 1065 1047 1081 1081
rect 991 1009 1081 1047
rect 1139 1081 1229 1097
rect 1139 1047 1155 1081
rect 1213 1047 1229 1081
rect 1139 1009 1229 1047
rect 1287 1081 1377 1097
rect 1287 1047 1303 1081
rect 1361 1047 1377 1081
rect 1287 1009 1377 1047
rect 1435 1081 1525 1097
rect 1435 1047 1451 1081
rect 1509 1047 1525 1081
rect 1435 1009 1525 1047
rect 1583 1081 1673 1097
rect 1583 1047 1599 1081
rect 1657 1047 1673 1081
rect 1583 1009 1673 1047
rect 1731 1081 1821 1097
rect 1731 1047 1747 1081
rect 1805 1047 1821 1081
rect 1731 1009 1821 1047
rect 1879 1081 1969 1097
rect 1879 1047 1895 1081
rect 1953 1047 1969 1081
rect 1879 1009 1969 1047
rect 2027 1081 2117 1097
rect 2027 1047 2043 1081
rect 2101 1047 2117 1081
rect 2027 1009 2117 1047
rect 2175 1081 2265 1097
rect 2175 1047 2191 1081
rect 2249 1047 2265 1081
rect 2175 1009 2265 1047
rect 2323 1081 2413 1097
rect 2323 1047 2339 1081
rect 2397 1047 2413 1081
rect 2323 1009 2413 1047
rect 2471 1081 2561 1097
rect 2471 1047 2487 1081
rect 2545 1047 2561 1081
rect 2471 1009 2561 1047
rect 2619 1081 2709 1097
rect 2619 1047 2635 1081
rect 2693 1047 2709 1081
rect 2619 1009 2709 1047
rect 2767 1081 2857 1097
rect 2767 1047 2783 1081
rect 2841 1047 2857 1081
rect 2767 1009 2857 1047
rect 2915 1081 3005 1097
rect 2915 1047 2931 1081
rect 2989 1047 3005 1081
rect 2915 1009 3005 1047
rect 3063 1081 3153 1097
rect 3063 1047 3079 1081
rect 3137 1047 3153 1081
rect 3063 1009 3153 1047
rect 3211 1081 3301 1097
rect 3211 1047 3227 1081
rect 3285 1047 3301 1081
rect 3211 1009 3301 1047
rect 3359 1081 3449 1097
rect 3359 1047 3375 1081
rect 3433 1047 3449 1081
rect 3359 1009 3449 1047
rect 3507 1081 3597 1097
rect 3507 1047 3523 1081
rect 3581 1047 3597 1081
rect 3507 1009 3597 1047
rect 3655 1081 3745 1097
rect 3655 1047 3671 1081
rect 3729 1047 3745 1081
rect 3655 1009 3745 1047
rect 3803 1081 3893 1097
rect 3803 1047 3819 1081
rect 3877 1047 3893 1081
rect 3803 1009 3893 1047
rect 3951 1081 4041 1097
rect 3951 1047 3967 1081
rect 4025 1047 4041 1081
rect 3951 1009 4041 1047
rect 4099 1081 4189 1097
rect 4099 1047 4115 1081
rect 4173 1047 4189 1081
rect 4099 1009 4189 1047
rect 4247 1081 4337 1097
rect 4247 1047 4263 1081
rect 4321 1047 4337 1081
rect 4247 1009 4337 1047
rect 4395 1081 4485 1097
rect 4395 1047 4411 1081
rect 4469 1047 4485 1081
rect 4395 1009 4485 1047
rect 4543 1081 4633 1097
rect 4543 1047 4559 1081
rect 4617 1047 4633 1081
rect 4543 1009 4633 1047
rect 4691 1081 4781 1097
rect 4691 1047 4707 1081
rect 4765 1047 4781 1081
rect 4691 1009 4781 1047
rect 4839 1081 4929 1097
rect 4839 1047 4855 1081
rect 4913 1047 4929 1081
rect 4839 1009 4929 1047
rect 4987 1081 5077 1097
rect 4987 1047 5003 1081
rect 5061 1047 5077 1081
rect 4987 1009 5077 1047
rect 5135 1081 5225 1097
rect 5135 1047 5151 1081
rect 5209 1047 5225 1081
rect 5135 1009 5225 1047
rect 5283 1081 5373 1097
rect 5283 1047 5299 1081
rect 5357 1047 5373 1081
rect 5283 1009 5373 1047
rect 5431 1081 5521 1097
rect 5431 1047 5447 1081
rect 5505 1047 5521 1081
rect 5431 1009 5521 1047
rect -5521 71 -5431 109
rect -5521 37 -5505 71
rect -5447 37 -5431 71
rect -5521 21 -5431 37
rect -5373 71 -5283 109
rect -5373 37 -5357 71
rect -5299 37 -5283 71
rect -5373 21 -5283 37
rect -5225 71 -5135 109
rect -5225 37 -5209 71
rect -5151 37 -5135 71
rect -5225 21 -5135 37
rect -5077 71 -4987 109
rect -5077 37 -5061 71
rect -5003 37 -4987 71
rect -5077 21 -4987 37
rect -4929 71 -4839 109
rect -4929 37 -4913 71
rect -4855 37 -4839 71
rect -4929 21 -4839 37
rect -4781 71 -4691 109
rect -4781 37 -4765 71
rect -4707 37 -4691 71
rect -4781 21 -4691 37
rect -4633 71 -4543 109
rect -4633 37 -4617 71
rect -4559 37 -4543 71
rect -4633 21 -4543 37
rect -4485 71 -4395 109
rect -4485 37 -4469 71
rect -4411 37 -4395 71
rect -4485 21 -4395 37
rect -4337 71 -4247 109
rect -4337 37 -4321 71
rect -4263 37 -4247 71
rect -4337 21 -4247 37
rect -4189 71 -4099 109
rect -4189 37 -4173 71
rect -4115 37 -4099 71
rect -4189 21 -4099 37
rect -4041 71 -3951 109
rect -4041 37 -4025 71
rect -3967 37 -3951 71
rect -4041 21 -3951 37
rect -3893 71 -3803 109
rect -3893 37 -3877 71
rect -3819 37 -3803 71
rect -3893 21 -3803 37
rect -3745 71 -3655 109
rect -3745 37 -3729 71
rect -3671 37 -3655 71
rect -3745 21 -3655 37
rect -3597 71 -3507 109
rect -3597 37 -3581 71
rect -3523 37 -3507 71
rect -3597 21 -3507 37
rect -3449 71 -3359 109
rect -3449 37 -3433 71
rect -3375 37 -3359 71
rect -3449 21 -3359 37
rect -3301 71 -3211 109
rect -3301 37 -3285 71
rect -3227 37 -3211 71
rect -3301 21 -3211 37
rect -3153 71 -3063 109
rect -3153 37 -3137 71
rect -3079 37 -3063 71
rect -3153 21 -3063 37
rect -3005 71 -2915 109
rect -3005 37 -2989 71
rect -2931 37 -2915 71
rect -3005 21 -2915 37
rect -2857 71 -2767 109
rect -2857 37 -2841 71
rect -2783 37 -2767 71
rect -2857 21 -2767 37
rect -2709 71 -2619 109
rect -2709 37 -2693 71
rect -2635 37 -2619 71
rect -2709 21 -2619 37
rect -2561 71 -2471 109
rect -2561 37 -2545 71
rect -2487 37 -2471 71
rect -2561 21 -2471 37
rect -2413 71 -2323 109
rect -2413 37 -2397 71
rect -2339 37 -2323 71
rect -2413 21 -2323 37
rect -2265 71 -2175 109
rect -2265 37 -2249 71
rect -2191 37 -2175 71
rect -2265 21 -2175 37
rect -2117 71 -2027 109
rect -2117 37 -2101 71
rect -2043 37 -2027 71
rect -2117 21 -2027 37
rect -1969 71 -1879 109
rect -1969 37 -1953 71
rect -1895 37 -1879 71
rect -1969 21 -1879 37
rect -1821 71 -1731 109
rect -1821 37 -1805 71
rect -1747 37 -1731 71
rect -1821 21 -1731 37
rect -1673 71 -1583 109
rect -1673 37 -1657 71
rect -1599 37 -1583 71
rect -1673 21 -1583 37
rect -1525 71 -1435 109
rect -1525 37 -1509 71
rect -1451 37 -1435 71
rect -1525 21 -1435 37
rect -1377 71 -1287 109
rect -1377 37 -1361 71
rect -1303 37 -1287 71
rect -1377 21 -1287 37
rect -1229 71 -1139 109
rect -1229 37 -1213 71
rect -1155 37 -1139 71
rect -1229 21 -1139 37
rect -1081 71 -991 109
rect -1081 37 -1065 71
rect -1007 37 -991 71
rect -1081 21 -991 37
rect -933 71 -843 109
rect -933 37 -917 71
rect -859 37 -843 71
rect -933 21 -843 37
rect -785 71 -695 109
rect -785 37 -769 71
rect -711 37 -695 71
rect -785 21 -695 37
rect -637 71 -547 109
rect -637 37 -621 71
rect -563 37 -547 71
rect -637 21 -547 37
rect -489 71 -399 109
rect -489 37 -473 71
rect -415 37 -399 71
rect -489 21 -399 37
rect -341 71 -251 109
rect -341 37 -325 71
rect -267 37 -251 71
rect -341 21 -251 37
rect -193 71 -103 109
rect -193 37 -177 71
rect -119 37 -103 71
rect -193 21 -103 37
rect -45 71 45 109
rect -45 37 -29 71
rect 29 37 45 71
rect -45 21 45 37
rect 103 71 193 109
rect 103 37 119 71
rect 177 37 193 71
rect 103 21 193 37
rect 251 71 341 109
rect 251 37 267 71
rect 325 37 341 71
rect 251 21 341 37
rect 399 71 489 109
rect 399 37 415 71
rect 473 37 489 71
rect 399 21 489 37
rect 547 71 637 109
rect 547 37 563 71
rect 621 37 637 71
rect 547 21 637 37
rect 695 71 785 109
rect 695 37 711 71
rect 769 37 785 71
rect 695 21 785 37
rect 843 71 933 109
rect 843 37 859 71
rect 917 37 933 71
rect 843 21 933 37
rect 991 71 1081 109
rect 991 37 1007 71
rect 1065 37 1081 71
rect 991 21 1081 37
rect 1139 71 1229 109
rect 1139 37 1155 71
rect 1213 37 1229 71
rect 1139 21 1229 37
rect 1287 71 1377 109
rect 1287 37 1303 71
rect 1361 37 1377 71
rect 1287 21 1377 37
rect 1435 71 1525 109
rect 1435 37 1451 71
rect 1509 37 1525 71
rect 1435 21 1525 37
rect 1583 71 1673 109
rect 1583 37 1599 71
rect 1657 37 1673 71
rect 1583 21 1673 37
rect 1731 71 1821 109
rect 1731 37 1747 71
rect 1805 37 1821 71
rect 1731 21 1821 37
rect 1879 71 1969 109
rect 1879 37 1895 71
rect 1953 37 1969 71
rect 1879 21 1969 37
rect 2027 71 2117 109
rect 2027 37 2043 71
rect 2101 37 2117 71
rect 2027 21 2117 37
rect 2175 71 2265 109
rect 2175 37 2191 71
rect 2249 37 2265 71
rect 2175 21 2265 37
rect 2323 71 2413 109
rect 2323 37 2339 71
rect 2397 37 2413 71
rect 2323 21 2413 37
rect 2471 71 2561 109
rect 2471 37 2487 71
rect 2545 37 2561 71
rect 2471 21 2561 37
rect 2619 71 2709 109
rect 2619 37 2635 71
rect 2693 37 2709 71
rect 2619 21 2709 37
rect 2767 71 2857 109
rect 2767 37 2783 71
rect 2841 37 2857 71
rect 2767 21 2857 37
rect 2915 71 3005 109
rect 2915 37 2931 71
rect 2989 37 3005 71
rect 2915 21 3005 37
rect 3063 71 3153 109
rect 3063 37 3079 71
rect 3137 37 3153 71
rect 3063 21 3153 37
rect 3211 71 3301 109
rect 3211 37 3227 71
rect 3285 37 3301 71
rect 3211 21 3301 37
rect 3359 71 3449 109
rect 3359 37 3375 71
rect 3433 37 3449 71
rect 3359 21 3449 37
rect 3507 71 3597 109
rect 3507 37 3523 71
rect 3581 37 3597 71
rect 3507 21 3597 37
rect 3655 71 3745 109
rect 3655 37 3671 71
rect 3729 37 3745 71
rect 3655 21 3745 37
rect 3803 71 3893 109
rect 3803 37 3819 71
rect 3877 37 3893 71
rect 3803 21 3893 37
rect 3951 71 4041 109
rect 3951 37 3967 71
rect 4025 37 4041 71
rect 3951 21 4041 37
rect 4099 71 4189 109
rect 4099 37 4115 71
rect 4173 37 4189 71
rect 4099 21 4189 37
rect 4247 71 4337 109
rect 4247 37 4263 71
rect 4321 37 4337 71
rect 4247 21 4337 37
rect 4395 71 4485 109
rect 4395 37 4411 71
rect 4469 37 4485 71
rect 4395 21 4485 37
rect 4543 71 4633 109
rect 4543 37 4559 71
rect 4617 37 4633 71
rect 4543 21 4633 37
rect 4691 71 4781 109
rect 4691 37 4707 71
rect 4765 37 4781 71
rect 4691 21 4781 37
rect 4839 71 4929 109
rect 4839 37 4855 71
rect 4913 37 4929 71
rect 4839 21 4929 37
rect 4987 71 5077 109
rect 4987 37 5003 71
rect 5061 37 5077 71
rect 4987 21 5077 37
rect 5135 71 5225 109
rect 5135 37 5151 71
rect 5209 37 5225 71
rect 5135 21 5225 37
rect 5283 71 5373 109
rect 5283 37 5299 71
rect 5357 37 5373 71
rect 5283 21 5373 37
rect 5431 71 5521 109
rect 5431 37 5447 71
rect 5505 37 5521 71
rect 5431 21 5521 37
rect -5521 -37 -5431 -21
rect -5521 -71 -5505 -37
rect -5447 -71 -5431 -37
rect -5521 -109 -5431 -71
rect -5373 -37 -5283 -21
rect -5373 -71 -5357 -37
rect -5299 -71 -5283 -37
rect -5373 -109 -5283 -71
rect -5225 -37 -5135 -21
rect -5225 -71 -5209 -37
rect -5151 -71 -5135 -37
rect -5225 -109 -5135 -71
rect -5077 -37 -4987 -21
rect -5077 -71 -5061 -37
rect -5003 -71 -4987 -37
rect -5077 -109 -4987 -71
rect -4929 -37 -4839 -21
rect -4929 -71 -4913 -37
rect -4855 -71 -4839 -37
rect -4929 -109 -4839 -71
rect -4781 -37 -4691 -21
rect -4781 -71 -4765 -37
rect -4707 -71 -4691 -37
rect -4781 -109 -4691 -71
rect -4633 -37 -4543 -21
rect -4633 -71 -4617 -37
rect -4559 -71 -4543 -37
rect -4633 -109 -4543 -71
rect -4485 -37 -4395 -21
rect -4485 -71 -4469 -37
rect -4411 -71 -4395 -37
rect -4485 -109 -4395 -71
rect -4337 -37 -4247 -21
rect -4337 -71 -4321 -37
rect -4263 -71 -4247 -37
rect -4337 -109 -4247 -71
rect -4189 -37 -4099 -21
rect -4189 -71 -4173 -37
rect -4115 -71 -4099 -37
rect -4189 -109 -4099 -71
rect -4041 -37 -3951 -21
rect -4041 -71 -4025 -37
rect -3967 -71 -3951 -37
rect -4041 -109 -3951 -71
rect -3893 -37 -3803 -21
rect -3893 -71 -3877 -37
rect -3819 -71 -3803 -37
rect -3893 -109 -3803 -71
rect -3745 -37 -3655 -21
rect -3745 -71 -3729 -37
rect -3671 -71 -3655 -37
rect -3745 -109 -3655 -71
rect -3597 -37 -3507 -21
rect -3597 -71 -3581 -37
rect -3523 -71 -3507 -37
rect -3597 -109 -3507 -71
rect -3449 -37 -3359 -21
rect -3449 -71 -3433 -37
rect -3375 -71 -3359 -37
rect -3449 -109 -3359 -71
rect -3301 -37 -3211 -21
rect -3301 -71 -3285 -37
rect -3227 -71 -3211 -37
rect -3301 -109 -3211 -71
rect -3153 -37 -3063 -21
rect -3153 -71 -3137 -37
rect -3079 -71 -3063 -37
rect -3153 -109 -3063 -71
rect -3005 -37 -2915 -21
rect -3005 -71 -2989 -37
rect -2931 -71 -2915 -37
rect -3005 -109 -2915 -71
rect -2857 -37 -2767 -21
rect -2857 -71 -2841 -37
rect -2783 -71 -2767 -37
rect -2857 -109 -2767 -71
rect -2709 -37 -2619 -21
rect -2709 -71 -2693 -37
rect -2635 -71 -2619 -37
rect -2709 -109 -2619 -71
rect -2561 -37 -2471 -21
rect -2561 -71 -2545 -37
rect -2487 -71 -2471 -37
rect -2561 -109 -2471 -71
rect -2413 -37 -2323 -21
rect -2413 -71 -2397 -37
rect -2339 -71 -2323 -37
rect -2413 -109 -2323 -71
rect -2265 -37 -2175 -21
rect -2265 -71 -2249 -37
rect -2191 -71 -2175 -37
rect -2265 -109 -2175 -71
rect -2117 -37 -2027 -21
rect -2117 -71 -2101 -37
rect -2043 -71 -2027 -37
rect -2117 -109 -2027 -71
rect -1969 -37 -1879 -21
rect -1969 -71 -1953 -37
rect -1895 -71 -1879 -37
rect -1969 -109 -1879 -71
rect -1821 -37 -1731 -21
rect -1821 -71 -1805 -37
rect -1747 -71 -1731 -37
rect -1821 -109 -1731 -71
rect -1673 -37 -1583 -21
rect -1673 -71 -1657 -37
rect -1599 -71 -1583 -37
rect -1673 -109 -1583 -71
rect -1525 -37 -1435 -21
rect -1525 -71 -1509 -37
rect -1451 -71 -1435 -37
rect -1525 -109 -1435 -71
rect -1377 -37 -1287 -21
rect -1377 -71 -1361 -37
rect -1303 -71 -1287 -37
rect -1377 -109 -1287 -71
rect -1229 -37 -1139 -21
rect -1229 -71 -1213 -37
rect -1155 -71 -1139 -37
rect -1229 -109 -1139 -71
rect -1081 -37 -991 -21
rect -1081 -71 -1065 -37
rect -1007 -71 -991 -37
rect -1081 -109 -991 -71
rect -933 -37 -843 -21
rect -933 -71 -917 -37
rect -859 -71 -843 -37
rect -933 -109 -843 -71
rect -785 -37 -695 -21
rect -785 -71 -769 -37
rect -711 -71 -695 -37
rect -785 -109 -695 -71
rect -637 -37 -547 -21
rect -637 -71 -621 -37
rect -563 -71 -547 -37
rect -637 -109 -547 -71
rect -489 -37 -399 -21
rect -489 -71 -473 -37
rect -415 -71 -399 -37
rect -489 -109 -399 -71
rect -341 -37 -251 -21
rect -341 -71 -325 -37
rect -267 -71 -251 -37
rect -341 -109 -251 -71
rect -193 -37 -103 -21
rect -193 -71 -177 -37
rect -119 -71 -103 -37
rect -193 -109 -103 -71
rect -45 -37 45 -21
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect -45 -109 45 -71
rect 103 -37 193 -21
rect 103 -71 119 -37
rect 177 -71 193 -37
rect 103 -109 193 -71
rect 251 -37 341 -21
rect 251 -71 267 -37
rect 325 -71 341 -37
rect 251 -109 341 -71
rect 399 -37 489 -21
rect 399 -71 415 -37
rect 473 -71 489 -37
rect 399 -109 489 -71
rect 547 -37 637 -21
rect 547 -71 563 -37
rect 621 -71 637 -37
rect 547 -109 637 -71
rect 695 -37 785 -21
rect 695 -71 711 -37
rect 769 -71 785 -37
rect 695 -109 785 -71
rect 843 -37 933 -21
rect 843 -71 859 -37
rect 917 -71 933 -37
rect 843 -109 933 -71
rect 991 -37 1081 -21
rect 991 -71 1007 -37
rect 1065 -71 1081 -37
rect 991 -109 1081 -71
rect 1139 -37 1229 -21
rect 1139 -71 1155 -37
rect 1213 -71 1229 -37
rect 1139 -109 1229 -71
rect 1287 -37 1377 -21
rect 1287 -71 1303 -37
rect 1361 -71 1377 -37
rect 1287 -109 1377 -71
rect 1435 -37 1525 -21
rect 1435 -71 1451 -37
rect 1509 -71 1525 -37
rect 1435 -109 1525 -71
rect 1583 -37 1673 -21
rect 1583 -71 1599 -37
rect 1657 -71 1673 -37
rect 1583 -109 1673 -71
rect 1731 -37 1821 -21
rect 1731 -71 1747 -37
rect 1805 -71 1821 -37
rect 1731 -109 1821 -71
rect 1879 -37 1969 -21
rect 1879 -71 1895 -37
rect 1953 -71 1969 -37
rect 1879 -109 1969 -71
rect 2027 -37 2117 -21
rect 2027 -71 2043 -37
rect 2101 -71 2117 -37
rect 2027 -109 2117 -71
rect 2175 -37 2265 -21
rect 2175 -71 2191 -37
rect 2249 -71 2265 -37
rect 2175 -109 2265 -71
rect 2323 -37 2413 -21
rect 2323 -71 2339 -37
rect 2397 -71 2413 -37
rect 2323 -109 2413 -71
rect 2471 -37 2561 -21
rect 2471 -71 2487 -37
rect 2545 -71 2561 -37
rect 2471 -109 2561 -71
rect 2619 -37 2709 -21
rect 2619 -71 2635 -37
rect 2693 -71 2709 -37
rect 2619 -109 2709 -71
rect 2767 -37 2857 -21
rect 2767 -71 2783 -37
rect 2841 -71 2857 -37
rect 2767 -109 2857 -71
rect 2915 -37 3005 -21
rect 2915 -71 2931 -37
rect 2989 -71 3005 -37
rect 2915 -109 3005 -71
rect 3063 -37 3153 -21
rect 3063 -71 3079 -37
rect 3137 -71 3153 -37
rect 3063 -109 3153 -71
rect 3211 -37 3301 -21
rect 3211 -71 3227 -37
rect 3285 -71 3301 -37
rect 3211 -109 3301 -71
rect 3359 -37 3449 -21
rect 3359 -71 3375 -37
rect 3433 -71 3449 -37
rect 3359 -109 3449 -71
rect 3507 -37 3597 -21
rect 3507 -71 3523 -37
rect 3581 -71 3597 -37
rect 3507 -109 3597 -71
rect 3655 -37 3745 -21
rect 3655 -71 3671 -37
rect 3729 -71 3745 -37
rect 3655 -109 3745 -71
rect 3803 -37 3893 -21
rect 3803 -71 3819 -37
rect 3877 -71 3893 -37
rect 3803 -109 3893 -71
rect 3951 -37 4041 -21
rect 3951 -71 3967 -37
rect 4025 -71 4041 -37
rect 3951 -109 4041 -71
rect 4099 -37 4189 -21
rect 4099 -71 4115 -37
rect 4173 -71 4189 -37
rect 4099 -109 4189 -71
rect 4247 -37 4337 -21
rect 4247 -71 4263 -37
rect 4321 -71 4337 -37
rect 4247 -109 4337 -71
rect 4395 -37 4485 -21
rect 4395 -71 4411 -37
rect 4469 -71 4485 -37
rect 4395 -109 4485 -71
rect 4543 -37 4633 -21
rect 4543 -71 4559 -37
rect 4617 -71 4633 -37
rect 4543 -109 4633 -71
rect 4691 -37 4781 -21
rect 4691 -71 4707 -37
rect 4765 -71 4781 -37
rect 4691 -109 4781 -71
rect 4839 -37 4929 -21
rect 4839 -71 4855 -37
rect 4913 -71 4929 -37
rect 4839 -109 4929 -71
rect 4987 -37 5077 -21
rect 4987 -71 5003 -37
rect 5061 -71 5077 -37
rect 4987 -109 5077 -71
rect 5135 -37 5225 -21
rect 5135 -71 5151 -37
rect 5209 -71 5225 -37
rect 5135 -109 5225 -71
rect 5283 -37 5373 -21
rect 5283 -71 5299 -37
rect 5357 -71 5373 -37
rect 5283 -109 5373 -71
rect 5431 -37 5521 -21
rect 5431 -71 5447 -37
rect 5505 -71 5521 -37
rect 5431 -109 5521 -71
rect -5521 -1047 -5431 -1009
rect -5521 -1081 -5505 -1047
rect -5447 -1081 -5431 -1047
rect -5521 -1097 -5431 -1081
rect -5373 -1047 -5283 -1009
rect -5373 -1081 -5357 -1047
rect -5299 -1081 -5283 -1047
rect -5373 -1097 -5283 -1081
rect -5225 -1047 -5135 -1009
rect -5225 -1081 -5209 -1047
rect -5151 -1081 -5135 -1047
rect -5225 -1097 -5135 -1081
rect -5077 -1047 -4987 -1009
rect -5077 -1081 -5061 -1047
rect -5003 -1081 -4987 -1047
rect -5077 -1097 -4987 -1081
rect -4929 -1047 -4839 -1009
rect -4929 -1081 -4913 -1047
rect -4855 -1081 -4839 -1047
rect -4929 -1097 -4839 -1081
rect -4781 -1047 -4691 -1009
rect -4781 -1081 -4765 -1047
rect -4707 -1081 -4691 -1047
rect -4781 -1097 -4691 -1081
rect -4633 -1047 -4543 -1009
rect -4633 -1081 -4617 -1047
rect -4559 -1081 -4543 -1047
rect -4633 -1097 -4543 -1081
rect -4485 -1047 -4395 -1009
rect -4485 -1081 -4469 -1047
rect -4411 -1081 -4395 -1047
rect -4485 -1097 -4395 -1081
rect -4337 -1047 -4247 -1009
rect -4337 -1081 -4321 -1047
rect -4263 -1081 -4247 -1047
rect -4337 -1097 -4247 -1081
rect -4189 -1047 -4099 -1009
rect -4189 -1081 -4173 -1047
rect -4115 -1081 -4099 -1047
rect -4189 -1097 -4099 -1081
rect -4041 -1047 -3951 -1009
rect -4041 -1081 -4025 -1047
rect -3967 -1081 -3951 -1047
rect -4041 -1097 -3951 -1081
rect -3893 -1047 -3803 -1009
rect -3893 -1081 -3877 -1047
rect -3819 -1081 -3803 -1047
rect -3893 -1097 -3803 -1081
rect -3745 -1047 -3655 -1009
rect -3745 -1081 -3729 -1047
rect -3671 -1081 -3655 -1047
rect -3745 -1097 -3655 -1081
rect -3597 -1047 -3507 -1009
rect -3597 -1081 -3581 -1047
rect -3523 -1081 -3507 -1047
rect -3597 -1097 -3507 -1081
rect -3449 -1047 -3359 -1009
rect -3449 -1081 -3433 -1047
rect -3375 -1081 -3359 -1047
rect -3449 -1097 -3359 -1081
rect -3301 -1047 -3211 -1009
rect -3301 -1081 -3285 -1047
rect -3227 -1081 -3211 -1047
rect -3301 -1097 -3211 -1081
rect -3153 -1047 -3063 -1009
rect -3153 -1081 -3137 -1047
rect -3079 -1081 -3063 -1047
rect -3153 -1097 -3063 -1081
rect -3005 -1047 -2915 -1009
rect -3005 -1081 -2989 -1047
rect -2931 -1081 -2915 -1047
rect -3005 -1097 -2915 -1081
rect -2857 -1047 -2767 -1009
rect -2857 -1081 -2841 -1047
rect -2783 -1081 -2767 -1047
rect -2857 -1097 -2767 -1081
rect -2709 -1047 -2619 -1009
rect -2709 -1081 -2693 -1047
rect -2635 -1081 -2619 -1047
rect -2709 -1097 -2619 -1081
rect -2561 -1047 -2471 -1009
rect -2561 -1081 -2545 -1047
rect -2487 -1081 -2471 -1047
rect -2561 -1097 -2471 -1081
rect -2413 -1047 -2323 -1009
rect -2413 -1081 -2397 -1047
rect -2339 -1081 -2323 -1047
rect -2413 -1097 -2323 -1081
rect -2265 -1047 -2175 -1009
rect -2265 -1081 -2249 -1047
rect -2191 -1081 -2175 -1047
rect -2265 -1097 -2175 -1081
rect -2117 -1047 -2027 -1009
rect -2117 -1081 -2101 -1047
rect -2043 -1081 -2027 -1047
rect -2117 -1097 -2027 -1081
rect -1969 -1047 -1879 -1009
rect -1969 -1081 -1953 -1047
rect -1895 -1081 -1879 -1047
rect -1969 -1097 -1879 -1081
rect -1821 -1047 -1731 -1009
rect -1821 -1081 -1805 -1047
rect -1747 -1081 -1731 -1047
rect -1821 -1097 -1731 -1081
rect -1673 -1047 -1583 -1009
rect -1673 -1081 -1657 -1047
rect -1599 -1081 -1583 -1047
rect -1673 -1097 -1583 -1081
rect -1525 -1047 -1435 -1009
rect -1525 -1081 -1509 -1047
rect -1451 -1081 -1435 -1047
rect -1525 -1097 -1435 -1081
rect -1377 -1047 -1287 -1009
rect -1377 -1081 -1361 -1047
rect -1303 -1081 -1287 -1047
rect -1377 -1097 -1287 -1081
rect -1229 -1047 -1139 -1009
rect -1229 -1081 -1213 -1047
rect -1155 -1081 -1139 -1047
rect -1229 -1097 -1139 -1081
rect -1081 -1047 -991 -1009
rect -1081 -1081 -1065 -1047
rect -1007 -1081 -991 -1047
rect -1081 -1097 -991 -1081
rect -933 -1047 -843 -1009
rect -933 -1081 -917 -1047
rect -859 -1081 -843 -1047
rect -933 -1097 -843 -1081
rect -785 -1047 -695 -1009
rect -785 -1081 -769 -1047
rect -711 -1081 -695 -1047
rect -785 -1097 -695 -1081
rect -637 -1047 -547 -1009
rect -637 -1081 -621 -1047
rect -563 -1081 -547 -1047
rect -637 -1097 -547 -1081
rect -489 -1047 -399 -1009
rect -489 -1081 -473 -1047
rect -415 -1081 -399 -1047
rect -489 -1097 -399 -1081
rect -341 -1047 -251 -1009
rect -341 -1081 -325 -1047
rect -267 -1081 -251 -1047
rect -341 -1097 -251 -1081
rect -193 -1047 -103 -1009
rect -193 -1081 -177 -1047
rect -119 -1081 -103 -1047
rect -193 -1097 -103 -1081
rect -45 -1047 45 -1009
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect -45 -1097 45 -1081
rect 103 -1047 193 -1009
rect 103 -1081 119 -1047
rect 177 -1081 193 -1047
rect 103 -1097 193 -1081
rect 251 -1047 341 -1009
rect 251 -1081 267 -1047
rect 325 -1081 341 -1047
rect 251 -1097 341 -1081
rect 399 -1047 489 -1009
rect 399 -1081 415 -1047
rect 473 -1081 489 -1047
rect 399 -1097 489 -1081
rect 547 -1047 637 -1009
rect 547 -1081 563 -1047
rect 621 -1081 637 -1047
rect 547 -1097 637 -1081
rect 695 -1047 785 -1009
rect 695 -1081 711 -1047
rect 769 -1081 785 -1047
rect 695 -1097 785 -1081
rect 843 -1047 933 -1009
rect 843 -1081 859 -1047
rect 917 -1081 933 -1047
rect 843 -1097 933 -1081
rect 991 -1047 1081 -1009
rect 991 -1081 1007 -1047
rect 1065 -1081 1081 -1047
rect 991 -1097 1081 -1081
rect 1139 -1047 1229 -1009
rect 1139 -1081 1155 -1047
rect 1213 -1081 1229 -1047
rect 1139 -1097 1229 -1081
rect 1287 -1047 1377 -1009
rect 1287 -1081 1303 -1047
rect 1361 -1081 1377 -1047
rect 1287 -1097 1377 -1081
rect 1435 -1047 1525 -1009
rect 1435 -1081 1451 -1047
rect 1509 -1081 1525 -1047
rect 1435 -1097 1525 -1081
rect 1583 -1047 1673 -1009
rect 1583 -1081 1599 -1047
rect 1657 -1081 1673 -1047
rect 1583 -1097 1673 -1081
rect 1731 -1047 1821 -1009
rect 1731 -1081 1747 -1047
rect 1805 -1081 1821 -1047
rect 1731 -1097 1821 -1081
rect 1879 -1047 1969 -1009
rect 1879 -1081 1895 -1047
rect 1953 -1081 1969 -1047
rect 1879 -1097 1969 -1081
rect 2027 -1047 2117 -1009
rect 2027 -1081 2043 -1047
rect 2101 -1081 2117 -1047
rect 2027 -1097 2117 -1081
rect 2175 -1047 2265 -1009
rect 2175 -1081 2191 -1047
rect 2249 -1081 2265 -1047
rect 2175 -1097 2265 -1081
rect 2323 -1047 2413 -1009
rect 2323 -1081 2339 -1047
rect 2397 -1081 2413 -1047
rect 2323 -1097 2413 -1081
rect 2471 -1047 2561 -1009
rect 2471 -1081 2487 -1047
rect 2545 -1081 2561 -1047
rect 2471 -1097 2561 -1081
rect 2619 -1047 2709 -1009
rect 2619 -1081 2635 -1047
rect 2693 -1081 2709 -1047
rect 2619 -1097 2709 -1081
rect 2767 -1047 2857 -1009
rect 2767 -1081 2783 -1047
rect 2841 -1081 2857 -1047
rect 2767 -1097 2857 -1081
rect 2915 -1047 3005 -1009
rect 2915 -1081 2931 -1047
rect 2989 -1081 3005 -1047
rect 2915 -1097 3005 -1081
rect 3063 -1047 3153 -1009
rect 3063 -1081 3079 -1047
rect 3137 -1081 3153 -1047
rect 3063 -1097 3153 -1081
rect 3211 -1047 3301 -1009
rect 3211 -1081 3227 -1047
rect 3285 -1081 3301 -1047
rect 3211 -1097 3301 -1081
rect 3359 -1047 3449 -1009
rect 3359 -1081 3375 -1047
rect 3433 -1081 3449 -1047
rect 3359 -1097 3449 -1081
rect 3507 -1047 3597 -1009
rect 3507 -1081 3523 -1047
rect 3581 -1081 3597 -1047
rect 3507 -1097 3597 -1081
rect 3655 -1047 3745 -1009
rect 3655 -1081 3671 -1047
rect 3729 -1081 3745 -1047
rect 3655 -1097 3745 -1081
rect 3803 -1047 3893 -1009
rect 3803 -1081 3819 -1047
rect 3877 -1081 3893 -1047
rect 3803 -1097 3893 -1081
rect 3951 -1047 4041 -1009
rect 3951 -1081 3967 -1047
rect 4025 -1081 4041 -1047
rect 3951 -1097 4041 -1081
rect 4099 -1047 4189 -1009
rect 4099 -1081 4115 -1047
rect 4173 -1081 4189 -1047
rect 4099 -1097 4189 -1081
rect 4247 -1047 4337 -1009
rect 4247 -1081 4263 -1047
rect 4321 -1081 4337 -1047
rect 4247 -1097 4337 -1081
rect 4395 -1047 4485 -1009
rect 4395 -1081 4411 -1047
rect 4469 -1081 4485 -1047
rect 4395 -1097 4485 -1081
rect 4543 -1047 4633 -1009
rect 4543 -1081 4559 -1047
rect 4617 -1081 4633 -1047
rect 4543 -1097 4633 -1081
rect 4691 -1047 4781 -1009
rect 4691 -1081 4707 -1047
rect 4765 -1081 4781 -1047
rect 4691 -1097 4781 -1081
rect 4839 -1047 4929 -1009
rect 4839 -1081 4855 -1047
rect 4913 -1081 4929 -1047
rect 4839 -1097 4929 -1081
rect 4987 -1047 5077 -1009
rect 4987 -1081 5003 -1047
rect 5061 -1081 5077 -1047
rect 4987 -1097 5077 -1081
rect 5135 -1047 5225 -1009
rect 5135 -1081 5151 -1047
rect 5209 -1081 5225 -1047
rect 5135 -1097 5225 -1081
rect 5283 -1047 5373 -1009
rect 5283 -1081 5299 -1047
rect 5357 -1081 5373 -1047
rect 5283 -1097 5373 -1081
rect 5431 -1047 5521 -1009
rect 5431 -1081 5447 -1047
rect 5505 -1081 5521 -1047
rect 5431 -1097 5521 -1081
<< polycont >>
rect -5505 1047 -5447 1081
rect -5357 1047 -5299 1081
rect -5209 1047 -5151 1081
rect -5061 1047 -5003 1081
rect -4913 1047 -4855 1081
rect -4765 1047 -4707 1081
rect -4617 1047 -4559 1081
rect -4469 1047 -4411 1081
rect -4321 1047 -4263 1081
rect -4173 1047 -4115 1081
rect -4025 1047 -3967 1081
rect -3877 1047 -3819 1081
rect -3729 1047 -3671 1081
rect -3581 1047 -3523 1081
rect -3433 1047 -3375 1081
rect -3285 1047 -3227 1081
rect -3137 1047 -3079 1081
rect -2989 1047 -2931 1081
rect -2841 1047 -2783 1081
rect -2693 1047 -2635 1081
rect -2545 1047 -2487 1081
rect -2397 1047 -2339 1081
rect -2249 1047 -2191 1081
rect -2101 1047 -2043 1081
rect -1953 1047 -1895 1081
rect -1805 1047 -1747 1081
rect -1657 1047 -1599 1081
rect -1509 1047 -1451 1081
rect -1361 1047 -1303 1081
rect -1213 1047 -1155 1081
rect -1065 1047 -1007 1081
rect -917 1047 -859 1081
rect -769 1047 -711 1081
rect -621 1047 -563 1081
rect -473 1047 -415 1081
rect -325 1047 -267 1081
rect -177 1047 -119 1081
rect -29 1047 29 1081
rect 119 1047 177 1081
rect 267 1047 325 1081
rect 415 1047 473 1081
rect 563 1047 621 1081
rect 711 1047 769 1081
rect 859 1047 917 1081
rect 1007 1047 1065 1081
rect 1155 1047 1213 1081
rect 1303 1047 1361 1081
rect 1451 1047 1509 1081
rect 1599 1047 1657 1081
rect 1747 1047 1805 1081
rect 1895 1047 1953 1081
rect 2043 1047 2101 1081
rect 2191 1047 2249 1081
rect 2339 1047 2397 1081
rect 2487 1047 2545 1081
rect 2635 1047 2693 1081
rect 2783 1047 2841 1081
rect 2931 1047 2989 1081
rect 3079 1047 3137 1081
rect 3227 1047 3285 1081
rect 3375 1047 3433 1081
rect 3523 1047 3581 1081
rect 3671 1047 3729 1081
rect 3819 1047 3877 1081
rect 3967 1047 4025 1081
rect 4115 1047 4173 1081
rect 4263 1047 4321 1081
rect 4411 1047 4469 1081
rect 4559 1047 4617 1081
rect 4707 1047 4765 1081
rect 4855 1047 4913 1081
rect 5003 1047 5061 1081
rect 5151 1047 5209 1081
rect 5299 1047 5357 1081
rect 5447 1047 5505 1081
rect -5505 37 -5447 71
rect -5357 37 -5299 71
rect -5209 37 -5151 71
rect -5061 37 -5003 71
rect -4913 37 -4855 71
rect -4765 37 -4707 71
rect -4617 37 -4559 71
rect -4469 37 -4411 71
rect -4321 37 -4263 71
rect -4173 37 -4115 71
rect -4025 37 -3967 71
rect -3877 37 -3819 71
rect -3729 37 -3671 71
rect -3581 37 -3523 71
rect -3433 37 -3375 71
rect -3285 37 -3227 71
rect -3137 37 -3079 71
rect -2989 37 -2931 71
rect -2841 37 -2783 71
rect -2693 37 -2635 71
rect -2545 37 -2487 71
rect -2397 37 -2339 71
rect -2249 37 -2191 71
rect -2101 37 -2043 71
rect -1953 37 -1895 71
rect -1805 37 -1747 71
rect -1657 37 -1599 71
rect -1509 37 -1451 71
rect -1361 37 -1303 71
rect -1213 37 -1155 71
rect -1065 37 -1007 71
rect -917 37 -859 71
rect -769 37 -711 71
rect -621 37 -563 71
rect -473 37 -415 71
rect -325 37 -267 71
rect -177 37 -119 71
rect -29 37 29 71
rect 119 37 177 71
rect 267 37 325 71
rect 415 37 473 71
rect 563 37 621 71
rect 711 37 769 71
rect 859 37 917 71
rect 1007 37 1065 71
rect 1155 37 1213 71
rect 1303 37 1361 71
rect 1451 37 1509 71
rect 1599 37 1657 71
rect 1747 37 1805 71
rect 1895 37 1953 71
rect 2043 37 2101 71
rect 2191 37 2249 71
rect 2339 37 2397 71
rect 2487 37 2545 71
rect 2635 37 2693 71
rect 2783 37 2841 71
rect 2931 37 2989 71
rect 3079 37 3137 71
rect 3227 37 3285 71
rect 3375 37 3433 71
rect 3523 37 3581 71
rect 3671 37 3729 71
rect 3819 37 3877 71
rect 3967 37 4025 71
rect 4115 37 4173 71
rect 4263 37 4321 71
rect 4411 37 4469 71
rect 4559 37 4617 71
rect 4707 37 4765 71
rect 4855 37 4913 71
rect 5003 37 5061 71
rect 5151 37 5209 71
rect 5299 37 5357 71
rect 5447 37 5505 71
rect -5505 -71 -5447 -37
rect -5357 -71 -5299 -37
rect -5209 -71 -5151 -37
rect -5061 -71 -5003 -37
rect -4913 -71 -4855 -37
rect -4765 -71 -4707 -37
rect -4617 -71 -4559 -37
rect -4469 -71 -4411 -37
rect -4321 -71 -4263 -37
rect -4173 -71 -4115 -37
rect -4025 -71 -3967 -37
rect -3877 -71 -3819 -37
rect -3729 -71 -3671 -37
rect -3581 -71 -3523 -37
rect -3433 -71 -3375 -37
rect -3285 -71 -3227 -37
rect -3137 -71 -3079 -37
rect -2989 -71 -2931 -37
rect -2841 -71 -2783 -37
rect -2693 -71 -2635 -37
rect -2545 -71 -2487 -37
rect -2397 -71 -2339 -37
rect -2249 -71 -2191 -37
rect -2101 -71 -2043 -37
rect -1953 -71 -1895 -37
rect -1805 -71 -1747 -37
rect -1657 -71 -1599 -37
rect -1509 -71 -1451 -37
rect -1361 -71 -1303 -37
rect -1213 -71 -1155 -37
rect -1065 -71 -1007 -37
rect -917 -71 -859 -37
rect -769 -71 -711 -37
rect -621 -71 -563 -37
rect -473 -71 -415 -37
rect -325 -71 -267 -37
rect -177 -71 -119 -37
rect -29 -71 29 -37
rect 119 -71 177 -37
rect 267 -71 325 -37
rect 415 -71 473 -37
rect 563 -71 621 -37
rect 711 -71 769 -37
rect 859 -71 917 -37
rect 1007 -71 1065 -37
rect 1155 -71 1213 -37
rect 1303 -71 1361 -37
rect 1451 -71 1509 -37
rect 1599 -71 1657 -37
rect 1747 -71 1805 -37
rect 1895 -71 1953 -37
rect 2043 -71 2101 -37
rect 2191 -71 2249 -37
rect 2339 -71 2397 -37
rect 2487 -71 2545 -37
rect 2635 -71 2693 -37
rect 2783 -71 2841 -37
rect 2931 -71 2989 -37
rect 3079 -71 3137 -37
rect 3227 -71 3285 -37
rect 3375 -71 3433 -37
rect 3523 -71 3581 -37
rect 3671 -71 3729 -37
rect 3819 -71 3877 -37
rect 3967 -71 4025 -37
rect 4115 -71 4173 -37
rect 4263 -71 4321 -37
rect 4411 -71 4469 -37
rect 4559 -71 4617 -37
rect 4707 -71 4765 -37
rect 4855 -71 4913 -37
rect 5003 -71 5061 -37
rect 5151 -71 5209 -37
rect 5299 -71 5357 -37
rect 5447 -71 5505 -37
rect -5505 -1081 -5447 -1047
rect -5357 -1081 -5299 -1047
rect -5209 -1081 -5151 -1047
rect -5061 -1081 -5003 -1047
rect -4913 -1081 -4855 -1047
rect -4765 -1081 -4707 -1047
rect -4617 -1081 -4559 -1047
rect -4469 -1081 -4411 -1047
rect -4321 -1081 -4263 -1047
rect -4173 -1081 -4115 -1047
rect -4025 -1081 -3967 -1047
rect -3877 -1081 -3819 -1047
rect -3729 -1081 -3671 -1047
rect -3581 -1081 -3523 -1047
rect -3433 -1081 -3375 -1047
rect -3285 -1081 -3227 -1047
rect -3137 -1081 -3079 -1047
rect -2989 -1081 -2931 -1047
rect -2841 -1081 -2783 -1047
rect -2693 -1081 -2635 -1047
rect -2545 -1081 -2487 -1047
rect -2397 -1081 -2339 -1047
rect -2249 -1081 -2191 -1047
rect -2101 -1081 -2043 -1047
rect -1953 -1081 -1895 -1047
rect -1805 -1081 -1747 -1047
rect -1657 -1081 -1599 -1047
rect -1509 -1081 -1451 -1047
rect -1361 -1081 -1303 -1047
rect -1213 -1081 -1155 -1047
rect -1065 -1081 -1007 -1047
rect -917 -1081 -859 -1047
rect -769 -1081 -711 -1047
rect -621 -1081 -563 -1047
rect -473 -1081 -415 -1047
rect -325 -1081 -267 -1047
rect -177 -1081 -119 -1047
rect -29 -1081 29 -1047
rect 119 -1081 177 -1047
rect 267 -1081 325 -1047
rect 415 -1081 473 -1047
rect 563 -1081 621 -1047
rect 711 -1081 769 -1047
rect 859 -1081 917 -1047
rect 1007 -1081 1065 -1047
rect 1155 -1081 1213 -1047
rect 1303 -1081 1361 -1047
rect 1451 -1081 1509 -1047
rect 1599 -1081 1657 -1047
rect 1747 -1081 1805 -1047
rect 1895 -1081 1953 -1047
rect 2043 -1081 2101 -1047
rect 2191 -1081 2249 -1047
rect 2339 -1081 2397 -1047
rect 2487 -1081 2545 -1047
rect 2635 -1081 2693 -1047
rect 2783 -1081 2841 -1047
rect 2931 -1081 2989 -1047
rect 3079 -1081 3137 -1047
rect 3227 -1081 3285 -1047
rect 3375 -1081 3433 -1047
rect 3523 -1081 3581 -1047
rect 3671 -1081 3729 -1047
rect 3819 -1081 3877 -1047
rect 3967 -1081 4025 -1047
rect 4115 -1081 4173 -1047
rect 4263 -1081 4321 -1047
rect 4411 -1081 4469 -1047
rect 4559 -1081 4617 -1047
rect 4707 -1081 4765 -1047
rect 4855 -1081 4913 -1047
rect 5003 -1081 5061 -1047
rect 5151 -1081 5209 -1047
rect 5299 -1081 5357 -1047
rect 5447 -1081 5505 -1047
<< locali >>
rect -5681 1149 -5585 1183
rect 5585 1149 5681 1183
rect -5681 1087 -5647 1149
rect 5647 1087 5681 1149
rect -5521 1047 -5505 1081
rect -5447 1047 -5431 1081
rect -5373 1047 -5357 1081
rect -5299 1047 -5283 1081
rect -5225 1047 -5209 1081
rect -5151 1047 -5135 1081
rect -5077 1047 -5061 1081
rect -5003 1047 -4987 1081
rect -4929 1047 -4913 1081
rect -4855 1047 -4839 1081
rect -4781 1047 -4765 1081
rect -4707 1047 -4691 1081
rect -4633 1047 -4617 1081
rect -4559 1047 -4543 1081
rect -4485 1047 -4469 1081
rect -4411 1047 -4395 1081
rect -4337 1047 -4321 1081
rect -4263 1047 -4247 1081
rect -4189 1047 -4173 1081
rect -4115 1047 -4099 1081
rect -4041 1047 -4025 1081
rect -3967 1047 -3951 1081
rect -3893 1047 -3877 1081
rect -3819 1047 -3803 1081
rect -3745 1047 -3729 1081
rect -3671 1047 -3655 1081
rect -3597 1047 -3581 1081
rect -3523 1047 -3507 1081
rect -3449 1047 -3433 1081
rect -3375 1047 -3359 1081
rect -3301 1047 -3285 1081
rect -3227 1047 -3211 1081
rect -3153 1047 -3137 1081
rect -3079 1047 -3063 1081
rect -3005 1047 -2989 1081
rect -2931 1047 -2915 1081
rect -2857 1047 -2841 1081
rect -2783 1047 -2767 1081
rect -2709 1047 -2693 1081
rect -2635 1047 -2619 1081
rect -2561 1047 -2545 1081
rect -2487 1047 -2471 1081
rect -2413 1047 -2397 1081
rect -2339 1047 -2323 1081
rect -2265 1047 -2249 1081
rect -2191 1047 -2175 1081
rect -2117 1047 -2101 1081
rect -2043 1047 -2027 1081
rect -1969 1047 -1953 1081
rect -1895 1047 -1879 1081
rect -1821 1047 -1805 1081
rect -1747 1047 -1731 1081
rect -1673 1047 -1657 1081
rect -1599 1047 -1583 1081
rect -1525 1047 -1509 1081
rect -1451 1047 -1435 1081
rect -1377 1047 -1361 1081
rect -1303 1047 -1287 1081
rect -1229 1047 -1213 1081
rect -1155 1047 -1139 1081
rect -1081 1047 -1065 1081
rect -1007 1047 -991 1081
rect -933 1047 -917 1081
rect -859 1047 -843 1081
rect -785 1047 -769 1081
rect -711 1047 -695 1081
rect -637 1047 -621 1081
rect -563 1047 -547 1081
rect -489 1047 -473 1081
rect -415 1047 -399 1081
rect -341 1047 -325 1081
rect -267 1047 -251 1081
rect -193 1047 -177 1081
rect -119 1047 -103 1081
rect -45 1047 -29 1081
rect 29 1047 45 1081
rect 103 1047 119 1081
rect 177 1047 193 1081
rect 251 1047 267 1081
rect 325 1047 341 1081
rect 399 1047 415 1081
rect 473 1047 489 1081
rect 547 1047 563 1081
rect 621 1047 637 1081
rect 695 1047 711 1081
rect 769 1047 785 1081
rect 843 1047 859 1081
rect 917 1047 933 1081
rect 991 1047 1007 1081
rect 1065 1047 1081 1081
rect 1139 1047 1155 1081
rect 1213 1047 1229 1081
rect 1287 1047 1303 1081
rect 1361 1047 1377 1081
rect 1435 1047 1451 1081
rect 1509 1047 1525 1081
rect 1583 1047 1599 1081
rect 1657 1047 1673 1081
rect 1731 1047 1747 1081
rect 1805 1047 1821 1081
rect 1879 1047 1895 1081
rect 1953 1047 1969 1081
rect 2027 1047 2043 1081
rect 2101 1047 2117 1081
rect 2175 1047 2191 1081
rect 2249 1047 2265 1081
rect 2323 1047 2339 1081
rect 2397 1047 2413 1081
rect 2471 1047 2487 1081
rect 2545 1047 2561 1081
rect 2619 1047 2635 1081
rect 2693 1047 2709 1081
rect 2767 1047 2783 1081
rect 2841 1047 2857 1081
rect 2915 1047 2931 1081
rect 2989 1047 3005 1081
rect 3063 1047 3079 1081
rect 3137 1047 3153 1081
rect 3211 1047 3227 1081
rect 3285 1047 3301 1081
rect 3359 1047 3375 1081
rect 3433 1047 3449 1081
rect 3507 1047 3523 1081
rect 3581 1047 3597 1081
rect 3655 1047 3671 1081
rect 3729 1047 3745 1081
rect 3803 1047 3819 1081
rect 3877 1047 3893 1081
rect 3951 1047 3967 1081
rect 4025 1047 4041 1081
rect 4099 1047 4115 1081
rect 4173 1047 4189 1081
rect 4247 1047 4263 1081
rect 4321 1047 4337 1081
rect 4395 1047 4411 1081
rect 4469 1047 4485 1081
rect 4543 1047 4559 1081
rect 4617 1047 4633 1081
rect 4691 1047 4707 1081
rect 4765 1047 4781 1081
rect 4839 1047 4855 1081
rect 4913 1047 4929 1081
rect 4987 1047 5003 1081
rect 5061 1047 5077 1081
rect 5135 1047 5151 1081
rect 5209 1047 5225 1081
rect 5283 1047 5299 1081
rect 5357 1047 5373 1081
rect 5431 1047 5447 1081
rect 5505 1047 5521 1081
rect -5567 997 -5533 1013
rect -5567 105 -5533 121
rect -5419 997 -5385 1013
rect -5419 105 -5385 121
rect -5271 997 -5237 1013
rect -5271 105 -5237 121
rect -5123 997 -5089 1013
rect -5123 105 -5089 121
rect -4975 997 -4941 1013
rect -4975 105 -4941 121
rect -4827 997 -4793 1013
rect -4827 105 -4793 121
rect -4679 997 -4645 1013
rect -4679 105 -4645 121
rect -4531 997 -4497 1013
rect -4531 105 -4497 121
rect -4383 997 -4349 1013
rect -4383 105 -4349 121
rect -4235 997 -4201 1013
rect -4235 105 -4201 121
rect -4087 997 -4053 1013
rect -4087 105 -4053 121
rect -3939 997 -3905 1013
rect -3939 105 -3905 121
rect -3791 997 -3757 1013
rect -3791 105 -3757 121
rect -3643 997 -3609 1013
rect -3643 105 -3609 121
rect -3495 997 -3461 1013
rect -3495 105 -3461 121
rect -3347 997 -3313 1013
rect -3347 105 -3313 121
rect -3199 997 -3165 1013
rect -3199 105 -3165 121
rect -3051 997 -3017 1013
rect -3051 105 -3017 121
rect -2903 997 -2869 1013
rect -2903 105 -2869 121
rect -2755 997 -2721 1013
rect -2755 105 -2721 121
rect -2607 997 -2573 1013
rect -2607 105 -2573 121
rect -2459 997 -2425 1013
rect -2459 105 -2425 121
rect -2311 997 -2277 1013
rect -2311 105 -2277 121
rect -2163 997 -2129 1013
rect -2163 105 -2129 121
rect -2015 997 -1981 1013
rect -2015 105 -1981 121
rect -1867 997 -1833 1013
rect -1867 105 -1833 121
rect -1719 997 -1685 1013
rect -1719 105 -1685 121
rect -1571 997 -1537 1013
rect -1571 105 -1537 121
rect -1423 997 -1389 1013
rect -1423 105 -1389 121
rect -1275 997 -1241 1013
rect -1275 105 -1241 121
rect -1127 997 -1093 1013
rect -1127 105 -1093 121
rect -979 997 -945 1013
rect -979 105 -945 121
rect -831 997 -797 1013
rect -831 105 -797 121
rect -683 997 -649 1013
rect -683 105 -649 121
rect -535 997 -501 1013
rect -535 105 -501 121
rect -387 997 -353 1013
rect -387 105 -353 121
rect -239 997 -205 1013
rect -239 105 -205 121
rect -91 997 -57 1013
rect -91 105 -57 121
rect 57 997 91 1013
rect 57 105 91 121
rect 205 997 239 1013
rect 205 105 239 121
rect 353 997 387 1013
rect 353 105 387 121
rect 501 997 535 1013
rect 501 105 535 121
rect 649 997 683 1013
rect 649 105 683 121
rect 797 997 831 1013
rect 797 105 831 121
rect 945 997 979 1013
rect 945 105 979 121
rect 1093 997 1127 1013
rect 1093 105 1127 121
rect 1241 997 1275 1013
rect 1241 105 1275 121
rect 1389 997 1423 1013
rect 1389 105 1423 121
rect 1537 997 1571 1013
rect 1537 105 1571 121
rect 1685 997 1719 1013
rect 1685 105 1719 121
rect 1833 997 1867 1013
rect 1833 105 1867 121
rect 1981 997 2015 1013
rect 1981 105 2015 121
rect 2129 997 2163 1013
rect 2129 105 2163 121
rect 2277 997 2311 1013
rect 2277 105 2311 121
rect 2425 997 2459 1013
rect 2425 105 2459 121
rect 2573 997 2607 1013
rect 2573 105 2607 121
rect 2721 997 2755 1013
rect 2721 105 2755 121
rect 2869 997 2903 1013
rect 2869 105 2903 121
rect 3017 997 3051 1013
rect 3017 105 3051 121
rect 3165 997 3199 1013
rect 3165 105 3199 121
rect 3313 997 3347 1013
rect 3313 105 3347 121
rect 3461 997 3495 1013
rect 3461 105 3495 121
rect 3609 997 3643 1013
rect 3609 105 3643 121
rect 3757 997 3791 1013
rect 3757 105 3791 121
rect 3905 997 3939 1013
rect 3905 105 3939 121
rect 4053 997 4087 1013
rect 4053 105 4087 121
rect 4201 997 4235 1013
rect 4201 105 4235 121
rect 4349 997 4383 1013
rect 4349 105 4383 121
rect 4497 997 4531 1013
rect 4497 105 4531 121
rect 4645 997 4679 1013
rect 4645 105 4679 121
rect 4793 997 4827 1013
rect 4793 105 4827 121
rect 4941 997 4975 1013
rect 4941 105 4975 121
rect 5089 997 5123 1013
rect 5089 105 5123 121
rect 5237 997 5271 1013
rect 5237 105 5271 121
rect 5385 997 5419 1013
rect 5385 105 5419 121
rect 5533 997 5567 1013
rect 5533 105 5567 121
rect -5521 37 -5505 71
rect -5447 37 -5431 71
rect -5373 37 -5357 71
rect -5299 37 -5283 71
rect -5225 37 -5209 71
rect -5151 37 -5135 71
rect -5077 37 -5061 71
rect -5003 37 -4987 71
rect -4929 37 -4913 71
rect -4855 37 -4839 71
rect -4781 37 -4765 71
rect -4707 37 -4691 71
rect -4633 37 -4617 71
rect -4559 37 -4543 71
rect -4485 37 -4469 71
rect -4411 37 -4395 71
rect -4337 37 -4321 71
rect -4263 37 -4247 71
rect -4189 37 -4173 71
rect -4115 37 -4099 71
rect -4041 37 -4025 71
rect -3967 37 -3951 71
rect -3893 37 -3877 71
rect -3819 37 -3803 71
rect -3745 37 -3729 71
rect -3671 37 -3655 71
rect -3597 37 -3581 71
rect -3523 37 -3507 71
rect -3449 37 -3433 71
rect -3375 37 -3359 71
rect -3301 37 -3285 71
rect -3227 37 -3211 71
rect -3153 37 -3137 71
rect -3079 37 -3063 71
rect -3005 37 -2989 71
rect -2931 37 -2915 71
rect -2857 37 -2841 71
rect -2783 37 -2767 71
rect -2709 37 -2693 71
rect -2635 37 -2619 71
rect -2561 37 -2545 71
rect -2487 37 -2471 71
rect -2413 37 -2397 71
rect -2339 37 -2323 71
rect -2265 37 -2249 71
rect -2191 37 -2175 71
rect -2117 37 -2101 71
rect -2043 37 -2027 71
rect -1969 37 -1953 71
rect -1895 37 -1879 71
rect -1821 37 -1805 71
rect -1747 37 -1731 71
rect -1673 37 -1657 71
rect -1599 37 -1583 71
rect -1525 37 -1509 71
rect -1451 37 -1435 71
rect -1377 37 -1361 71
rect -1303 37 -1287 71
rect -1229 37 -1213 71
rect -1155 37 -1139 71
rect -1081 37 -1065 71
rect -1007 37 -991 71
rect -933 37 -917 71
rect -859 37 -843 71
rect -785 37 -769 71
rect -711 37 -695 71
rect -637 37 -621 71
rect -563 37 -547 71
rect -489 37 -473 71
rect -415 37 -399 71
rect -341 37 -325 71
rect -267 37 -251 71
rect -193 37 -177 71
rect -119 37 -103 71
rect -45 37 -29 71
rect 29 37 45 71
rect 103 37 119 71
rect 177 37 193 71
rect 251 37 267 71
rect 325 37 341 71
rect 399 37 415 71
rect 473 37 489 71
rect 547 37 563 71
rect 621 37 637 71
rect 695 37 711 71
rect 769 37 785 71
rect 843 37 859 71
rect 917 37 933 71
rect 991 37 1007 71
rect 1065 37 1081 71
rect 1139 37 1155 71
rect 1213 37 1229 71
rect 1287 37 1303 71
rect 1361 37 1377 71
rect 1435 37 1451 71
rect 1509 37 1525 71
rect 1583 37 1599 71
rect 1657 37 1673 71
rect 1731 37 1747 71
rect 1805 37 1821 71
rect 1879 37 1895 71
rect 1953 37 1969 71
rect 2027 37 2043 71
rect 2101 37 2117 71
rect 2175 37 2191 71
rect 2249 37 2265 71
rect 2323 37 2339 71
rect 2397 37 2413 71
rect 2471 37 2487 71
rect 2545 37 2561 71
rect 2619 37 2635 71
rect 2693 37 2709 71
rect 2767 37 2783 71
rect 2841 37 2857 71
rect 2915 37 2931 71
rect 2989 37 3005 71
rect 3063 37 3079 71
rect 3137 37 3153 71
rect 3211 37 3227 71
rect 3285 37 3301 71
rect 3359 37 3375 71
rect 3433 37 3449 71
rect 3507 37 3523 71
rect 3581 37 3597 71
rect 3655 37 3671 71
rect 3729 37 3745 71
rect 3803 37 3819 71
rect 3877 37 3893 71
rect 3951 37 3967 71
rect 4025 37 4041 71
rect 4099 37 4115 71
rect 4173 37 4189 71
rect 4247 37 4263 71
rect 4321 37 4337 71
rect 4395 37 4411 71
rect 4469 37 4485 71
rect 4543 37 4559 71
rect 4617 37 4633 71
rect 4691 37 4707 71
rect 4765 37 4781 71
rect 4839 37 4855 71
rect 4913 37 4929 71
rect 4987 37 5003 71
rect 5061 37 5077 71
rect 5135 37 5151 71
rect 5209 37 5225 71
rect 5283 37 5299 71
rect 5357 37 5373 71
rect 5431 37 5447 71
rect 5505 37 5521 71
rect -5521 -71 -5505 -37
rect -5447 -71 -5431 -37
rect -5373 -71 -5357 -37
rect -5299 -71 -5283 -37
rect -5225 -71 -5209 -37
rect -5151 -71 -5135 -37
rect -5077 -71 -5061 -37
rect -5003 -71 -4987 -37
rect -4929 -71 -4913 -37
rect -4855 -71 -4839 -37
rect -4781 -71 -4765 -37
rect -4707 -71 -4691 -37
rect -4633 -71 -4617 -37
rect -4559 -71 -4543 -37
rect -4485 -71 -4469 -37
rect -4411 -71 -4395 -37
rect -4337 -71 -4321 -37
rect -4263 -71 -4247 -37
rect -4189 -71 -4173 -37
rect -4115 -71 -4099 -37
rect -4041 -71 -4025 -37
rect -3967 -71 -3951 -37
rect -3893 -71 -3877 -37
rect -3819 -71 -3803 -37
rect -3745 -71 -3729 -37
rect -3671 -71 -3655 -37
rect -3597 -71 -3581 -37
rect -3523 -71 -3507 -37
rect -3449 -71 -3433 -37
rect -3375 -71 -3359 -37
rect -3301 -71 -3285 -37
rect -3227 -71 -3211 -37
rect -3153 -71 -3137 -37
rect -3079 -71 -3063 -37
rect -3005 -71 -2989 -37
rect -2931 -71 -2915 -37
rect -2857 -71 -2841 -37
rect -2783 -71 -2767 -37
rect -2709 -71 -2693 -37
rect -2635 -71 -2619 -37
rect -2561 -71 -2545 -37
rect -2487 -71 -2471 -37
rect -2413 -71 -2397 -37
rect -2339 -71 -2323 -37
rect -2265 -71 -2249 -37
rect -2191 -71 -2175 -37
rect -2117 -71 -2101 -37
rect -2043 -71 -2027 -37
rect -1969 -71 -1953 -37
rect -1895 -71 -1879 -37
rect -1821 -71 -1805 -37
rect -1747 -71 -1731 -37
rect -1673 -71 -1657 -37
rect -1599 -71 -1583 -37
rect -1525 -71 -1509 -37
rect -1451 -71 -1435 -37
rect -1377 -71 -1361 -37
rect -1303 -71 -1287 -37
rect -1229 -71 -1213 -37
rect -1155 -71 -1139 -37
rect -1081 -71 -1065 -37
rect -1007 -71 -991 -37
rect -933 -71 -917 -37
rect -859 -71 -843 -37
rect -785 -71 -769 -37
rect -711 -71 -695 -37
rect -637 -71 -621 -37
rect -563 -71 -547 -37
rect -489 -71 -473 -37
rect -415 -71 -399 -37
rect -341 -71 -325 -37
rect -267 -71 -251 -37
rect -193 -71 -177 -37
rect -119 -71 -103 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 103 -71 119 -37
rect 177 -71 193 -37
rect 251 -71 267 -37
rect 325 -71 341 -37
rect 399 -71 415 -37
rect 473 -71 489 -37
rect 547 -71 563 -37
rect 621 -71 637 -37
rect 695 -71 711 -37
rect 769 -71 785 -37
rect 843 -71 859 -37
rect 917 -71 933 -37
rect 991 -71 1007 -37
rect 1065 -71 1081 -37
rect 1139 -71 1155 -37
rect 1213 -71 1229 -37
rect 1287 -71 1303 -37
rect 1361 -71 1377 -37
rect 1435 -71 1451 -37
rect 1509 -71 1525 -37
rect 1583 -71 1599 -37
rect 1657 -71 1673 -37
rect 1731 -71 1747 -37
rect 1805 -71 1821 -37
rect 1879 -71 1895 -37
rect 1953 -71 1969 -37
rect 2027 -71 2043 -37
rect 2101 -71 2117 -37
rect 2175 -71 2191 -37
rect 2249 -71 2265 -37
rect 2323 -71 2339 -37
rect 2397 -71 2413 -37
rect 2471 -71 2487 -37
rect 2545 -71 2561 -37
rect 2619 -71 2635 -37
rect 2693 -71 2709 -37
rect 2767 -71 2783 -37
rect 2841 -71 2857 -37
rect 2915 -71 2931 -37
rect 2989 -71 3005 -37
rect 3063 -71 3079 -37
rect 3137 -71 3153 -37
rect 3211 -71 3227 -37
rect 3285 -71 3301 -37
rect 3359 -71 3375 -37
rect 3433 -71 3449 -37
rect 3507 -71 3523 -37
rect 3581 -71 3597 -37
rect 3655 -71 3671 -37
rect 3729 -71 3745 -37
rect 3803 -71 3819 -37
rect 3877 -71 3893 -37
rect 3951 -71 3967 -37
rect 4025 -71 4041 -37
rect 4099 -71 4115 -37
rect 4173 -71 4189 -37
rect 4247 -71 4263 -37
rect 4321 -71 4337 -37
rect 4395 -71 4411 -37
rect 4469 -71 4485 -37
rect 4543 -71 4559 -37
rect 4617 -71 4633 -37
rect 4691 -71 4707 -37
rect 4765 -71 4781 -37
rect 4839 -71 4855 -37
rect 4913 -71 4929 -37
rect 4987 -71 5003 -37
rect 5061 -71 5077 -37
rect 5135 -71 5151 -37
rect 5209 -71 5225 -37
rect 5283 -71 5299 -37
rect 5357 -71 5373 -37
rect 5431 -71 5447 -37
rect 5505 -71 5521 -37
rect -5567 -121 -5533 -105
rect -5567 -1013 -5533 -997
rect -5419 -121 -5385 -105
rect -5419 -1013 -5385 -997
rect -5271 -121 -5237 -105
rect -5271 -1013 -5237 -997
rect -5123 -121 -5089 -105
rect -5123 -1013 -5089 -997
rect -4975 -121 -4941 -105
rect -4975 -1013 -4941 -997
rect -4827 -121 -4793 -105
rect -4827 -1013 -4793 -997
rect -4679 -121 -4645 -105
rect -4679 -1013 -4645 -997
rect -4531 -121 -4497 -105
rect -4531 -1013 -4497 -997
rect -4383 -121 -4349 -105
rect -4383 -1013 -4349 -997
rect -4235 -121 -4201 -105
rect -4235 -1013 -4201 -997
rect -4087 -121 -4053 -105
rect -4087 -1013 -4053 -997
rect -3939 -121 -3905 -105
rect -3939 -1013 -3905 -997
rect -3791 -121 -3757 -105
rect -3791 -1013 -3757 -997
rect -3643 -121 -3609 -105
rect -3643 -1013 -3609 -997
rect -3495 -121 -3461 -105
rect -3495 -1013 -3461 -997
rect -3347 -121 -3313 -105
rect -3347 -1013 -3313 -997
rect -3199 -121 -3165 -105
rect -3199 -1013 -3165 -997
rect -3051 -121 -3017 -105
rect -3051 -1013 -3017 -997
rect -2903 -121 -2869 -105
rect -2903 -1013 -2869 -997
rect -2755 -121 -2721 -105
rect -2755 -1013 -2721 -997
rect -2607 -121 -2573 -105
rect -2607 -1013 -2573 -997
rect -2459 -121 -2425 -105
rect -2459 -1013 -2425 -997
rect -2311 -121 -2277 -105
rect -2311 -1013 -2277 -997
rect -2163 -121 -2129 -105
rect -2163 -1013 -2129 -997
rect -2015 -121 -1981 -105
rect -2015 -1013 -1981 -997
rect -1867 -121 -1833 -105
rect -1867 -1013 -1833 -997
rect -1719 -121 -1685 -105
rect -1719 -1013 -1685 -997
rect -1571 -121 -1537 -105
rect -1571 -1013 -1537 -997
rect -1423 -121 -1389 -105
rect -1423 -1013 -1389 -997
rect -1275 -121 -1241 -105
rect -1275 -1013 -1241 -997
rect -1127 -121 -1093 -105
rect -1127 -1013 -1093 -997
rect -979 -121 -945 -105
rect -979 -1013 -945 -997
rect -831 -121 -797 -105
rect -831 -1013 -797 -997
rect -683 -121 -649 -105
rect -683 -1013 -649 -997
rect -535 -121 -501 -105
rect -535 -1013 -501 -997
rect -387 -121 -353 -105
rect -387 -1013 -353 -997
rect -239 -121 -205 -105
rect -239 -1013 -205 -997
rect -91 -121 -57 -105
rect -91 -1013 -57 -997
rect 57 -121 91 -105
rect 57 -1013 91 -997
rect 205 -121 239 -105
rect 205 -1013 239 -997
rect 353 -121 387 -105
rect 353 -1013 387 -997
rect 501 -121 535 -105
rect 501 -1013 535 -997
rect 649 -121 683 -105
rect 649 -1013 683 -997
rect 797 -121 831 -105
rect 797 -1013 831 -997
rect 945 -121 979 -105
rect 945 -1013 979 -997
rect 1093 -121 1127 -105
rect 1093 -1013 1127 -997
rect 1241 -121 1275 -105
rect 1241 -1013 1275 -997
rect 1389 -121 1423 -105
rect 1389 -1013 1423 -997
rect 1537 -121 1571 -105
rect 1537 -1013 1571 -997
rect 1685 -121 1719 -105
rect 1685 -1013 1719 -997
rect 1833 -121 1867 -105
rect 1833 -1013 1867 -997
rect 1981 -121 2015 -105
rect 1981 -1013 2015 -997
rect 2129 -121 2163 -105
rect 2129 -1013 2163 -997
rect 2277 -121 2311 -105
rect 2277 -1013 2311 -997
rect 2425 -121 2459 -105
rect 2425 -1013 2459 -997
rect 2573 -121 2607 -105
rect 2573 -1013 2607 -997
rect 2721 -121 2755 -105
rect 2721 -1013 2755 -997
rect 2869 -121 2903 -105
rect 2869 -1013 2903 -997
rect 3017 -121 3051 -105
rect 3017 -1013 3051 -997
rect 3165 -121 3199 -105
rect 3165 -1013 3199 -997
rect 3313 -121 3347 -105
rect 3313 -1013 3347 -997
rect 3461 -121 3495 -105
rect 3461 -1013 3495 -997
rect 3609 -121 3643 -105
rect 3609 -1013 3643 -997
rect 3757 -121 3791 -105
rect 3757 -1013 3791 -997
rect 3905 -121 3939 -105
rect 3905 -1013 3939 -997
rect 4053 -121 4087 -105
rect 4053 -1013 4087 -997
rect 4201 -121 4235 -105
rect 4201 -1013 4235 -997
rect 4349 -121 4383 -105
rect 4349 -1013 4383 -997
rect 4497 -121 4531 -105
rect 4497 -1013 4531 -997
rect 4645 -121 4679 -105
rect 4645 -1013 4679 -997
rect 4793 -121 4827 -105
rect 4793 -1013 4827 -997
rect 4941 -121 4975 -105
rect 4941 -1013 4975 -997
rect 5089 -121 5123 -105
rect 5089 -1013 5123 -997
rect 5237 -121 5271 -105
rect 5237 -1013 5271 -997
rect 5385 -121 5419 -105
rect 5385 -1013 5419 -997
rect 5533 -121 5567 -105
rect 5533 -1013 5567 -997
rect -5521 -1081 -5505 -1047
rect -5447 -1081 -5431 -1047
rect -5373 -1081 -5357 -1047
rect -5299 -1081 -5283 -1047
rect -5225 -1081 -5209 -1047
rect -5151 -1081 -5135 -1047
rect -5077 -1081 -5061 -1047
rect -5003 -1081 -4987 -1047
rect -4929 -1081 -4913 -1047
rect -4855 -1081 -4839 -1047
rect -4781 -1081 -4765 -1047
rect -4707 -1081 -4691 -1047
rect -4633 -1081 -4617 -1047
rect -4559 -1081 -4543 -1047
rect -4485 -1081 -4469 -1047
rect -4411 -1081 -4395 -1047
rect -4337 -1081 -4321 -1047
rect -4263 -1081 -4247 -1047
rect -4189 -1081 -4173 -1047
rect -4115 -1081 -4099 -1047
rect -4041 -1081 -4025 -1047
rect -3967 -1081 -3951 -1047
rect -3893 -1081 -3877 -1047
rect -3819 -1081 -3803 -1047
rect -3745 -1081 -3729 -1047
rect -3671 -1081 -3655 -1047
rect -3597 -1081 -3581 -1047
rect -3523 -1081 -3507 -1047
rect -3449 -1081 -3433 -1047
rect -3375 -1081 -3359 -1047
rect -3301 -1081 -3285 -1047
rect -3227 -1081 -3211 -1047
rect -3153 -1081 -3137 -1047
rect -3079 -1081 -3063 -1047
rect -3005 -1081 -2989 -1047
rect -2931 -1081 -2915 -1047
rect -2857 -1081 -2841 -1047
rect -2783 -1081 -2767 -1047
rect -2709 -1081 -2693 -1047
rect -2635 -1081 -2619 -1047
rect -2561 -1081 -2545 -1047
rect -2487 -1081 -2471 -1047
rect -2413 -1081 -2397 -1047
rect -2339 -1081 -2323 -1047
rect -2265 -1081 -2249 -1047
rect -2191 -1081 -2175 -1047
rect -2117 -1081 -2101 -1047
rect -2043 -1081 -2027 -1047
rect -1969 -1081 -1953 -1047
rect -1895 -1081 -1879 -1047
rect -1821 -1081 -1805 -1047
rect -1747 -1081 -1731 -1047
rect -1673 -1081 -1657 -1047
rect -1599 -1081 -1583 -1047
rect -1525 -1081 -1509 -1047
rect -1451 -1081 -1435 -1047
rect -1377 -1081 -1361 -1047
rect -1303 -1081 -1287 -1047
rect -1229 -1081 -1213 -1047
rect -1155 -1081 -1139 -1047
rect -1081 -1081 -1065 -1047
rect -1007 -1081 -991 -1047
rect -933 -1081 -917 -1047
rect -859 -1081 -843 -1047
rect -785 -1081 -769 -1047
rect -711 -1081 -695 -1047
rect -637 -1081 -621 -1047
rect -563 -1081 -547 -1047
rect -489 -1081 -473 -1047
rect -415 -1081 -399 -1047
rect -341 -1081 -325 -1047
rect -267 -1081 -251 -1047
rect -193 -1081 -177 -1047
rect -119 -1081 -103 -1047
rect -45 -1081 -29 -1047
rect 29 -1081 45 -1047
rect 103 -1081 119 -1047
rect 177 -1081 193 -1047
rect 251 -1081 267 -1047
rect 325 -1081 341 -1047
rect 399 -1081 415 -1047
rect 473 -1081 489 -1047
rect 547 -1081 563 -1047
rect 621 -1081 637 -1047
rect 695 -1081 711 -1047
rect 769 -1081 785 -1047
rect 843 -1081 859 -1047
rect 917 -1081 933 -1047
rect 991 -1081 1007 -1047
rect 1065 -1081 1081 -1047
rect 1139 -1081 1155 -1047
rect 1213 -1081 1229 -1047
rect 1287 -1081 1303 -1047
rect 1361 -1081 1377 -1047
rect 1435 -1081 1451 -1047
rect 1509 -1081 1525 -1047
rect 1583 -1081 1599 -1047
rect 1657 -1081 1673 -1047
rect 1731 -1081 1747 -1047
rect 1805 -1081 1821 -1047
rect 1879 -1081 1895 -1047
rect 1953 -1081 1969 -1047
rect 2027 -1081 2043 -1047
rect 2101 -1081 2117 -1047
rect 2175 -1081 2191 -1047
rect 2249 -1081 2265 -1047
rect 2323 -1081 2339 -1047
rect 2397 -1081 2413 -1047
rect 2471 -1081 2487 -1047
rect 2545 -1081 2561 -1047
rect 2619 -1081 2635 -1047
rect 2693 -1081 2709 -1047
rect 2767 -1081 2783 -1047
rect 2841 -1081 2857 -1047
rect 2915 -1081 2931 -1047
rect 2989 -1081 3005 -1047
rect 3063 -1081 3079 -1047
rect 3137 -1081 3153 -1047
rect 3211 -1081 3227 -1047
rect 3285 -1081 3301 -1047
rect 3359 -1081 3375 -1047
rect 3433 -1081 3449 -1047
rect 3507 -1081 3523 -1047
rect 3581 -1081 3597 -1047
rect 3655 -1081 3671 -1047
rect 3729 -1081 3745 -1047
rect 3803 -1081 3819 -1047
rect 3877 -1081 3893 -1047
rect 3951 -1081 3967 -1047
rect 4025 -1081 4041 -1047
rect 4099 -1081 4115 -1047
rect 4173 -1081 4189 -1047
rect 4247 -1081 4263 -1047
rect 4321 -1081 4337 -1047
rect 4395 -1081 4411 -1047
rect 4469 -1081 4485 -1047
rect 4543 -1081 4559 -1047
rect 4617 -1081 4633 -1047
rect 4691 -1081 4707 -1047
rect 4765 -1081 4781 -1047
rect 4839 -1081 4855 -1047
rect 4913 -1081 4929 -1047
rect 4987 -1081 5003 -1047
rect 5061 -1081 5077 -1047
rect 5135 -1081 5151 -1047
rect 5209 -1081 5225 -1047
rect 5283 -1081 5299 -1047
rect 5357 -1081 5373 -1047
rect 5431 -1081 5447 -1047
rect 5505 -1081 5521 -1047
rect -5681 -1149 -5647 -1087
rect 5647 -1149 5681 -1087
rect -5681 -1183 -5585 -1149
rect 5585 -1183 5681 -1149
<< viali >>
rect -5505 1047 -5447 1081
rect -5357 1047 -5299 1081
rect -5209 1047 -5151 1081
rect -5061 1047 -5003 1081
rect -4913 1047 -4855 1081
rect -4765 1047 -4707 1081
rect -4617 1047 -4559 1081
rect -4469 1047 -4411 1081
rect -4321 1047 -4263 1081
rect -4173 1047 -4115 1081
rect -4025 1047 -3967 1081
rect -3877 1047 -3819 1081
rect -3729 1047 -3671 1081
rect -3581 1047 -3523 1081
rect -3433 1047 -3375 1081
rect -3285 1047 -3227 1081
rect -3137 1047 -3079 1081
rect -2989 1047 -2931 1081
rect -2841 1047 -2783 1081
rect -2693 1047 -2635 1081
rect -2545 1047 -2487 1081
rect -2397 1047 -2339 1081
rect -2249 1047 -2191 1081
rect -2101 1047 -2043 1081
rect -1953 1047 -1895 1081
rect -1805 1047 -1747 1081
rect -1657 1047 -1599 1081
rect -1509 1047 -1451 1081
rect -1361 1047 -1303 1081
rect -1213 1047 -1155 1081
rect -1065 1047 -1007 1081
rect -917 1047 -859 1081
rect -769 1047 -711 1081
rect -621 1047 -563 1081
rect -473 1047 -415 1081
rect -325 1047 -267 1081
rect -177 1047 -119 1081
rect -29 1047 29 1081
rect 119 1047 177 1081
rect 267 1047 325 1081
rect 415 1047 473 1081
rect 563 1047 621 1081
rect 711 1047 769 1081
rect 859 1047 917 1081
rect 1007 1047 1065 1081
rect 1155 1047 1213 1081
rect 1303 1047 1361 1081
rect 1451 1047 1509 1081
rect 1599 1047 1657 1081
rect 1747 1047 1805 1081
rect 1895 1047 1953 1081
rect 2043 1047 2101 1081
rect 2191 1047 2249 1081
rect 2339 1047 2397 1081
rect 2487 1047 2545 1081
rect 2635 1047 2693 1081
rect 2783 1047 2841 1081
rect 2931 1047 2989 1081
rect 3079 1047 3137 1081
rect 3227 1047 3285 1081
rect 3375 1047 3433 1081
rect 3523 1047 3581 1081
rect 3671 1047 3729 1081
rect 3819 1047 3877 1081
rect 3967 1047 4025 1081
rect 4115 1047 4173 1081
rect 4263 1047 4321 1081
rect 4411 1047 4469 1081
rect 4559 1047 4617 1081
rect 4707 1047 4765 1081
rect 4855 1047 4913 1081
rect 5003 1047 5061 1081
rect 5151 1047 5209 1081
rect 5299 1047 5357 1081
rect 5447 1047 5505 1081
rect -5567 121 -5533 997
rect -5419 121 -5385 997
rect -5271 121 -5237 997
rect -5123 121 -5089 997
rect -4975 121 -4941 997
rect -4827 121 -4793 997
rect -4679 121 -4645 997
rect -4531 121 -4497 997
rect -4383 121 -4349 997
rect -4235 121 -4201 997
rect -4087 121 -4053 997
rect -3939 121 -3905 997
rect -3791 121 -3757 997
rect -3643 121 -3609 997
rect -3495 121 -3461 997
rect -3347 121 -3313 997
rect -3199 121 -3165 997
rect -3051 121 -3017 997
rect -2903 121 -2869 997
rect -2755 121 -2721 997
rect -2607 121 -2573 997
rect -2459 121 -2425 997
rect -2311 121 -2277 997
rect -2163 121 -2129 997
rect -2015 121 -1981 997
rect -1867 121 -1833 997
rect -1719 121 -1685 997
rect -1571 121 -1537 997
rect -1423 121 -1389 997
rect -1275 121 -1241 997
rect -1127 121 -1093 997
rect -979 121 -945 997
rect -831 121 -797 997
rect -683 121 -649 997
rect -535 121 -501 997
rect -387 121 -353 997
rect -239 121 -205 997
rect -91 121 -57 997
rect 57 121 91 997
rect 205 121 239 997
rect 353 121 387 997
rect 501 121 535 997
rect 649 121 683 997
rect 797 121 831 997
rect 945 121 979 997
rect 1093 121 1127 997
rect 1241 121 1275 997
rect 1389 121 1423 997
rect 1537 121 1571 997
rect 1685 121 1719 997
rect 1833 121 1867 997
rect 1981 121 2015 997
rect 2129 121 2163 997
rect 2277 121 2311 997
rect 2425 121 2459 997
rect 2573 121 2607 997
rect 2721 121 2755 997
rect 2869 121 2903 997
rect 3017 121 3051 997
rect 3165 121 3199 997
rect 3313 121 3347 997
rect 3461 121 3495 997
rect 3609 121 3643 997
rect 3757 121 3791 997
rect 3905 121 3939 997
rect 4053 121 4087 997
rect 4201 121 4235 997
rect 4349 121 4383 997
rect 4497 121 4531 997
rect 4645 121 4679 997
rect 4793 121 4827 997
rect 4941 121 4975 997
rect 5089 121 5123 997
rect 5237 121 5271 997
rect 5385 121 5419 997
rect 5533 121 5567 997
rect -5505 37 -5447 71
rect -5357 37 -5299 71
rect -5209 37 -5151 71
rect -5061 37 -5003 71
rect -4913 37 -4855 71
rect -4765 37 -4707 71
rect -4617 37 -4559 71
rect -4469 37 -4411 71
rect -4321 37 -4263 71
rect -4173 37 -4115 71
rect -4025 37 -3967 71
rect -3877 37 -3819 71
rect -3729 37 -3671 71
rect -3581 37 -3523 71
rect -3433 37 -3375 71
rect -3285 37 -3227 71
rect -3137 37 -3079 71
rect -2989 37 -2931 71
rect -2841 37 -2783 71
rect -2693 37 -2635 71
rect -2545 37 -2487 71
rect -2397 37 -2339 71
rect -2249 37 -2191 71
rect -2101 37 -2043 71
rect -1953 37 -1895 71
rect -1805 37 -1747 71
rect -1657 37 -1599 71
rect -1509 37 -1451 71
rect -1361 37 -1303 71
rect -1213 37 -1155 71
rect -1065 37 -1007 71
rect -917 37 -859 71
rect -769 37 -711 71
rect -621 37 -563 71
rect -473 37 -415 71
rect -325 37 -267 71
rect -177 37 -119 71
rect -29 37 29 71
rect 119 37 177 71
rect 267 37 325 71
rect 415 37 473 71
rect 563 37 621 71
rect 711 37 769 71
rect 859 37 917 71
rect 1007 37 1065 71
rect 1155 37 1213 71
rect 1303 37 1361 71
rect 1451 37 1509 71
rect 1599 37 1657 71
rect 1747 37 1805 71
rect 1895 37 1953 71
rect 2043 37 2101 71
rect 2191 37 2249 71
rect 2339 37 2397 71
rect 2487 37 2545 71
rect 2635 37 2693 71
rect 2783 37 2841 71
rect 2931 37 2989 71
rect 3079 37 3137 71
rect 3227 37 3285 71
rect 3375 37 3433 71
rect 3523 37 3581 71
rect 3671 37 3729 71
rect 3819 37 3877 71
rect 3967 37 4025 71
rect 4115 37 4173 71
rect 4263 37 4321 71
rect 4411 37 4469 71
rect 4559 37 4617 71
rect 4707 37 4765 71
rect 4855 37 4913 71
rect 5003 37 5061 71
rect 5151 37 5209 71
rect 5299 37 5357 71
rect 5447 37 5505 71
rect -5505 -71 -5447 -37
rect -5357 -71 -5299 -37
rect -5209 -71 -5151 -37
rect -5061 -71 -5003 -37
rect -4913 -71 -4855 -37
rect -4765 -71 -4707 -37
rect -4617 -71 -4559 -37
rect -4469 -71 -4411 -37
rect -4321 -71 -4263 -37
rect -4173 -71 -4115 -37
rect -4025 -71 -3967 -37
rect -3877 -71 -3819 -37
rect -3729 -71 -3671 -37
rect -3581 -71 -3523 -37
rect -3433 -71 -3375 -37
rect -3285 -71 -3227 -37
rect -3137 -71 -3079 -37
rect -2989 -71 -2931 -37
rect -2841 -71 -2783 -37
rect -2693 -71 -2635 -37
rect -2545 -71 -2487 -37
rect -2397 -71 -2339 -37
rect -2249 -71 -2191 -37
rect -2101 -71 -2043 -37
rect -1953 -71 -1895 -37
rect -1805 -71 -1747 -37
rect -1657 -71 -1599 -37
rect -1509 -71 -1451 -37
rect -1361 -71 -1303 -37
rect -1213 -71 -1155 -37
rect -1065 -71 -1007 -37
rect -917 -71 -859 -37
rect -769 -71 -711 -37
rect -621 -71 -563 -37
rect -473 -71 -415 -37
rect -325 -71 -267 -37
rect -177 -71 -119 -37
rect -29 -71 29 -37
rect 119 -71 177 -37
rect 267 -71 325 -37
rect 415 -71 473 -37
rect 563 -71 621 -37
rect 711 -71 769 -37
rect 859 -71 917 -37
rect 1007 -71 1065 -37
rect 1155 -71 1213 -37
rect 1303 -71 1361 -37
rect 1451 -71 1509 -37
rect 1599 -71 1657 -37
rect 1747 -71 1805 -37
rect 1895 -71 1953 -37
rect 2043 -71 2101 -37
rect 2191 -71 2249 -37
rect 2339 -71 2397 -37
rect 2487 -71 2545 -37
rect 2635 -71 2693 -37
rect 2783 -71 2841 -37
rect 2931 -71 2989 -37
rect 3079 -71 3137 -37
rect 3227 -71 3285 -37
rect 3375 -71 3433 -37
rect 3523 -71 3581 -37
rect 3671 -71 3729 -37
rect 3819 -71 3877 -37
rect 3967 -71 4025 -37
rect 4115 -71 4173 -37
rect 4263 -71 4321 -37
rect 4411 -71 4469 -37
rect 4559 -71 4617 -37
rect 4707 -71 4765 -37
rect 4855 -71 4913 -37
rect 5003 -71 5061 -37
rect 5151 -71 5209 -37
rect 5299 -71 5357 -37
rect 5447 -71 5505 -37
rect -5567 -997 -5533 -121
rect -5419 -997 -5385 -121
rect -5271 -997 -5237 -121
rect -5123 -997 -5089 -121
rect -4975 -997 -4941 -121
rect -4827 -997 -4793 -121
rect -4679 -997 -4645 -121
rect -4531 -997 -4497 -121
rect -4383 -997 -4349 -121
rect -4235 -997 -4201 -121
rect -4087 -997 -4053 -121
rect -3939 -997 -3905 -121
rect -3791 -997 -3757 -121
rect -3643 -997 -3609 -121
rect -3495 -997 -3461 -121
rect -3347 -997 -3313 -121
rect -3199 -997 -3165 -121
rect -3051 -997 -3017 -121
rect -2903 -997 -2869 -121
rect -2755 -997 -2721 -121
rect -2607 -997 -2573 -121
rect -2459 -997 -2425 -121
rect -2311 -997 -2277 -121
rect -2163 -997 -2129 -121
rect -2015 -997 -1981 -121
rect -1867 -997 -1833 -121
rect -1719 -997 -1685 -121
rect -1571 -997 -1537 -121
rect -1423 -997 -1389 -121
rect -1275 -997 -1241 -121
rect -1127 -997 -1093 -121
rect -979 -997 -945 -121
rect -831 -997 -797 -121
rect -683 -997 -649 -121
rect -535 -997 -501 -121
rect -387 -997 -353 -121
rect -239 -997 -205 -121
rect -91 -997 -57 -121
rect 57 -997 91 -121
rect 205 -997 239 -121
rect 353 -997 387 -121
rect 501 -997 535 -121
rect 649 -997 683 -121
rect 797 -997 831 -121
rect 945 -997 979 -121
rect 1093 -997 1127 -121
rect 1241 -997 1275 -121
rect 1389 -997 1423 -121
rect 1537 -997 1571 -121
rect 1685 -997 1719 -121
rect 1833 -997 1867 -121
rect 1981 -997 2015 -121
rect 2129 -997 2163 -121
rect 2277 -997 2311 -121
rect 2425 -997 2459 -121
rect 2573 -997 2607 -121
rect 2721 -997 2755 -121
rect 2869 -997 2903 -121
rect 3017 -997 3051 -121
rect 3165 -997 3199 -121
rect 3313 -997 3347 -121
rect 3461 -997 3495 -121
rect 3609 -997 3643 -121
rect 3757 -997 3791 -121
rect 3905 -997 3939 -121
rect 4053 -997 4087 -121
rect 4201 -997 4235 -121
rect 4349 -997 4383 -121
rect 4497 -997 4531 -121
rect 4645 -997 4679 -121
rect 4793 -997 4827 -121
rect 4941 -997 4975 -121
rect 5089 -997 5123 -121
rect 5237 -997 5271 -121
rect 5385 -997 5419 -121
rect 5533 -997 5567 -121
rect -5505 -1081 -5447 -1047
rect -5357 -1081 -5299 -1047
rect -5209 -1081 -5151 -1047
rect -5061 -1081 -5003 -1047
rect -4913 -1081 -4855 -1047
rect -4765 -1081 -4707 -1047
rect -4617 -1081 -4559 -1047
rect -4469 -1081 -4411 -1047
rect -4321 -1081 -4263 -1047
rect -4173 -1081 -4115 -1047
rect -4025 -1081 -3967 -1047
rect -3877 -1081 -3819 -1047
rect -3729 -1081 -3671 -1047
rect -3581 -1081 -3523 -1047
rect -3433 -1081 -3375 -1047
rect -3285 -1081 -3227 -1047
rect -3137 -1081 -3079 -1047
rect -2989 -1081 -2931 -1047
rect -2841 -1081 -2783 -1047
rect -2693 -1081 -2635 -1047
rect -2545 -1081 -2487 -1047
rect -2397 -1081 -2339 -1047
rect -2249 -1081 -2191 -1047
rect -2101 -1081 -2043 -1047
rect -1953 -1081 -1895 -1047
rect -1805 -1081 -1747 -1047
rect -1657 -1081 -1599 -1047
rect -1509 -1081 -1451 -1047
rect -1361 -1081 -1303 -1047
rect -1213 -1081 -1155 -1047
rect -1065 -1081 -1007 -1047
rect -917 -1081 -859 -1047
rect -769 -1081 -711 -1047
rect -621 -1081 -563 -1047
rect -473 -1081 -415 -1047
rect -325 -1081 -267 -1047
rect -177 -1081 -119 -1047
rect -29 -1081 29 -1047
rect 119 -1081 177 -1047
rect 267 -1081 325 -1047
rect 415 -1081 473 -1047
rect 563 -1081 621 -1047
rect 711 -1081 769 -1047
rect 859 -1081 917 -1047
rect 1007 -1081 1065 -1047
rect 1155 -1081 1213 -1047
rect 1303 -1081 1361 -1047
rect 1451 -1081 1509 -1047
rect 1599 -1081 1657 -1047
rect 1747 -1081 1805 -1047
rect 1895 -1081 1953 -1047
rect 2043 -1081 2101 -1047
rect 2191 -1081 2249 -1047
rect 2339 -1081 2397 -1047
rect 2487 -1081 2545 -1047
rect 2635 -1081 2693 -1047
rect 2783 -1081 2841 -1047
rect 2931 -1081 2989 -1047
rect 3079 -1081 3137 -1047
rect 3227 -1081 3285 -1047
rect 3375 -1081 3433 -1047
rect 3523 -1081 3581 -1047
rect 3671 -1081 3729 -1047
rect 3819 -1081 3877 -1047
rect 3967 -1081 4025 -1047
rect 4115 -1081 4173 -1047
rect 4263 -1081 4321 -1047
rect 4411 -1081 4469 -1047
rect 4559 -1081 4617 -1047
rect 4707 -1081 4765 -1047
rect 4855 -1081 4913 -1047
rect 5003 -1081 5061 -1047
rect 5151 -1081 5209 -1047
rect 5299 -1081 5357 -1047
rect 5447 -1081 5505 -1047
<< metal1 >>
rect -5517 1081 -5435 1087
rect -5517 1047 -5505 1081
rect -5447 1047 -5435 1081
rect -5517 1041 -5435 1047
rect -5369 1081 -5287 1087
rect -5369 1047 -5357 1081
rect -5299 1047 -5287 1081
rect -5369 1041 -5287 1047
rect -5221 1081 -5139 1087
rect -5221 1047 -5209 1081
rect -5151 1047 -5139 1081
rect -5221 1041 -5139 1047
rect -5073 1081 -4991 1087
rect -5073 1047 -5061 1081
rect -5003 1047 -4991 1081
rect -5073 1041 -4991 1047
rect -4925 1081 -4843 1087
rect -4925 1047 -4913 1081
rect -4855 1047 -4843 1081
rect -4925 1041 -4843 1047
rect -4777 1081 -4695 1087
rect -4777 1047 -4765 1081
rect -4707 1047 -4695 1081
rect -4777 1041 -4695 1047
rect -4629 1081 -4547 1087
rect -4629 1047 -4617 1081
rect -4559 1047 -4547 1081
rect -4629 1041 -4547 1047
rect -4481 1081 -4399 1087
rect -4481 1047 -4469 1081
rect -4411 1047 -4399 1081
rect -4481 1041 -4399 1047
rect -4333 1081 -4251 1087
rect -4333 1047 -4321 1081
rect -4263 1047 -4251 1081
rect -4333 1041 -4251 1047
rect -4185 1081 -4103 1087
rect -4185 1047 -4173 1081
rect -4115 1047 -4103 1081
rect -4185 1041 -4103 1047
rect -4037 1081 -3955 1087
rect -4037 1047 -4025 1081
rect -3967 1047 -3955 1081
rect -4037 1041 -3955 1047
rect -3889 1081 -3807 1087
rect -3889 1047 -3877 1081
rect -3819 1047 -3807 1081
rect -3889 1041 -3807 1047
rect -3741 1081 -3659 1087
rect -3741 1047 -3729 1081
rect -3671 1047 -3659 1081
rect -3741 1041 -3659 1047
rect -3593 1081 -3511 1087
rect -3593 1047 -3581 1081
rect -3523 1047 -3511 1081
rect -3593 1041 -3511 1047
rect -3445 1081 -3363 1087
rect -3445 1047 -3433 1081
rect -3375 1047 -3363 1081
rect -3445 1041 -3363 1047
rect -3297 1081 -3215 1087
rect -3297 1047 -3285 1081
rect -3227 1047 -3215 1081
rect -3297 1041 -3215 1047
rect -3149 1081 -3067 1087
rect -3149 1047 -3137 1081
rect -3079 1047 -3067 1081
rect -3149 1041 -3067 1047
rect -3001 1081 -2919 1087
rect -3001 1047 -2989 1081
rect -2931 1047 -2919 1081
rect -3001 1041 -2919 1047
rect -2853 1081 -2771 1087
rect -2853 1047 -2841 1081
rect -2783 1047 -2771 1081
rect -2853 1041 -2771 1047
rect -2705 1081 -2623 1087
rect -2705 1047 -2693 1081
rect -2635 1047 -2623 1081
rect -2705 1041 -2623 1047
rect -2557 1081 -2475 1087
rect -2557 1047 -2545 1081
rect -2487 1047 -2475 1081
rect -2557 1041 -2475 1047
rect -2409 1081 -2327 1087
rect -2409 1047 -2397 1081
rect -2339 1047 -2327 1081
rect -2409 1041 -2327 1047
rect -2261 1081 -2179 1087
rect -2261 1047 -2249 1081
rect -2191 1047 -2179 1081
rect -2261 1041 -2179 1047
rect -2113 1081 -2031 1087
rect -2113 1047 -2101 1081
rect -2043 1047 -2031 1081
rect -2113 1041 -2031 1047
rect -1965 1081 -1883 1087
rect -1965 1047 -1953 1081
rect -1895 1047 -1883 1081
rect -1965 1041 -1883 1047
rect -1817 1081 -1735 1087
rect -1817 1047 -1805 1081
rect -1747 1047 -1735 1081
rect -1817 1041 -1735 1047
rect -1669 1081 -1587 1087
rect -1669 1047 -1657 1081
rect -1599 1047 -1587 1081
rect -1669 1041 -1587 1047
rect -1521 1081 -1439 1087
rect -1521 1047 -1509 1081
rect -1451 1047 -1439 1081
rect -1521 1041 -1439 1047
rect -1373 1081 -1291 1087
rect -1373 1047 -1361 1081
rect -1303 1047 -1291 1081
rect -1373 1041 -1291 1047
rect -1225 1081 -1143 1087
rect -1225 1047 -1213 1081
rect -1155 1047 -1143 1081
rect -1225 1041 -1143 1047
rect -1077 1081 -995 1087
rect -1077 1047 -1065 1081
rect -1007 1047 -995 1081
rect -1077 1041 -995 1047
rect -929 1081 -847 1087
rect -929 1047 -917 1081
rect -859 1047 -847 1081
rect -929 1041 -847 1047
rect -781 1081 -699 1087
rect -781 1047 -769 1081
rect -711 1047 -699 1081
rect -781 1041 -699 1047
rect -633 1081 -551 1087
rect -633 1047 -621 1081
rect -563 1047 -551 1081
rect -633 1041 -551 1047
rect -485 1081 -403 1087
rect -485 1047 -473 1081
rect -415 1047 -403 1081
rect -485 1041 -403 1047
rect -337 1081 -255 1087
rect -337 1047 -325 1081
rect -267 1047 -255 1081
rect -337 1041 -255 1047
rect -189 1081 -107 1087
rect -189 1047 -177 1081
rect -119 1047 -107 1081
rect -189 1041 -107 1047
rect -41 1081 41 1087
rect -41 1047 -29 1081
rect 29 1047 41 1081
rect -41 1041 41 1047
rect 107 1081 189 1087
rect 107 1047 119 1081
rect 177 1047 189 1081
rect 107 1041 189 1047
rect 255 1081 337 1087
rect 255 1047 267 1081
rect 325 1047 337 1081
rect 255 1041 337 1047
rect 403 1081 485 1087
rect 403 1047 415 1081
rect 473 1047 485 1081
rect 403 1041 485 1047
rect 551 1081 633 1087
rect 551 1047 563 1081
rect 621 1047 633 1081
rect 551 1041 633 1047
rect 699 1081 781 1087
rect 699 1047 711 1081
rect 769 1047 781 1081
rect 699 1041 781 1047
rect 847 1081 929 1087
rect 847 1047 859 1081
rect 917 1047 929 1081
rect 847 1041 929 1047
rect 995 1081 1077 1087
rect 995 1047 1007 1081
rect 1065 1047 1077 1081
rect 995 1041 1077 1047
rect 1143 1081 1225 1087
rect 1143 1047 1155 1081
rect 1213 1047 1225 1081
rect 1143 1041 1225 1047
rect 1291 1081 1373 1087
rect 1291 1047 1303 1081
rect 1361 1047 1373 1081
rect 1291 1041 1373 1047
rect 1439 1081 1521 1087
rect 1439 1047 1451 1081
rect 1509 1047 1521 1081
rect 1439 1041 1521 1047
rect 1587 1081 1669 1087
rect 1587 1047 1599 1081
rect 1657 1047 1669 1081
rect 1587 1041 1669 1047
rect 1735 1081 1817 1087
rect 1735 1047 1747 1081
rect 1805 1047 1817 1081
rect 1735 1041 1817 1047
rect 1883 1081 1965 1087
rect 1883 1047 1895 1081
rect 1953 1047 1965 1081
rect 1883 1041 1965 1047
rect 2031 1081 2113 1087
rect 2031 1047 2043 1081
rect 2101 1047 2113 1081
rect 2031 1041 2113 1047
rect 2179 1081 2261 1087
rect 2179 1047 2191 1081
rect 2249 1047 2261 1081
rect 2179 1041 2261 1047
rect 2327 1081 2409 1087
rect 2327 1047 2339 1081
rect 2397 1047 2409 1081
rect 2327 1041 2409 1047
rect 2475 1081 2557 1087
rect 2475 1047 2487 1081
rect 2545 1047 2557 1081
rect 2475 1041 2557 1047
rect 2623 1081 2705 1087
rect 2623 1047 2635 1081
rect 2693 1047 2705 1081
rect 2623 1041 2705 1047
rect 2771 1081 2853 1087
rect 2771 1047 2783 1081
rect 2841 1047 2853 1081
rect 2771 1041 2853 1047
rect 2919 1081 3001 1087
rect 2919 1047 2931 1081
rect 2989 1047 3001 1081
rect 2919 1041 3001 1047
rect 3067 1081 3149 1087
rect 3067 1047 3079 1081
rect 3137 1047 3149 1081
rect 3067 1041 3149 1047
rect 3215 1081 3297 1087
rect 3215 1047 3227 1081
rect 3285 1047 3297 1081
rect 3215 1041 3297 1047
rect 3363 1081 3445 1087
rect 3363 1047 3375 1081
rect 3433 1047 3445 1081
rect 3363 1041 3445 1047
rect 3511 1081 3593 1087
rect 3511 1047 3523 1081
rect 3581 1047 3593 1081
rect 3511 1041 3593 1047
rect 3659 1081 3741 1087
rect 3659 1047 3671 1081
rect 3729 1047 3741 1081
rect 3659 1041 3741 1047
rect 3807 1081 3889 1087
rect 3807 1047 3819 1081
rect 3877 1047 3889 1081
rect 3807 1041 3889 1047
rect 3955 1081 4037 1087
rect 3955 1047 3967 1081
rect 4025 1047 4037 1081
rect 3955 1041 4037 1047
rect 4103 1081 4185 1087
rect 4103 1047 4115 1081
rect 4173 1047 4185 1081
rect 4103 1041 4185 1047
rect 4251 1081 4333 1087
rect 4251 1047 4263 1081
rect 4321 1047 4333 1081
rect 4251 1041 4333 1047
rect 4399 1081 4481 1087
rect 4399 1047 4411 1081
rect 4469 1047 4481 1081
rect 4399 1041 4481 1047
rect 4547 1081 4629 1087
rect 4547 1047 4559 1081
rect 4617 1047 4629 1081
rect 4547 1041 4629 1047
rect 4695 1081 4777 1087
rect 4695 1047 4707 1081
rect 4765 1047 4777 1081
rect 4695 1041 4777 1047
rect 4843 1081 4925 1087
rect 4843 1047 4855 1081
rect 4913 1047 4925 1081
rect 4843 1041 4925 1047
rect 4991 1081 5073 1087
rect 4991 1047 5003 1081
rect 5061 1047 5073 1081
rect 4991 1041 5073 1047
rect 5139 1081 5221 1087
rect 5139 1047 5151 1081
rect 5209 1047 5221 1081
rect 5139 1041 5221 1047
rect 5287 1081 5369 1087
rect 5287 1047 5299 1081
rect 5357 1047 5369 1081
rect 5287 1041 5369 1047
rect 5435 1081 5517 1087
rect 5435 1047 5447 1081
rect 5505 1047 5517 1081
rect 5435 1041 5517 1047
rect -5573 997 -5527 1009
rect -5573 121 -5567 997
rect -5533 121 -5527 997
rect -5573 109 -5527 121
rect -5425 997 -5379 1009
rect -5425 121 -5419 997
rect -5385 121 -5379 997
rect -5425 109 -5379 121
rect -5277 997 -5231 1009
rect -5277 121 -5271 997
rect -5237 121 -5231 997
rect -5277 109 -5231 121
rect -5129 997 -5083 1009
rect -5129 121 -5123 997
rect -5089 121 -5083 997
rect -5129 109 -5083 121
rect -4981 997 -4935 1009
rect -4981 121 -4975 997
rect -4941 121 -4935 997
rect -4981 109 -4935 121
rect -4833 997 -4787 1009
rect -4833 121 -4827 997
rect -4793 121 -4787 997
rect -4833 109 -4787 121
rect -4685 997 -4639 1009
rect -4685 121 -4679 997
rect -4645 121 -4639 997
rect -4685 109 -4639 121
rect -4537 997 -4491 1009
rect -4537 121 -4531 997
rect -4497 121 -4491 997
rect -4537 109 -4491 121
rect -4389 997 -4343 1009
rect -4389 121 -4383 997
rect -4349 121 -4343 997
rect -4389 109 -4343 121
rect -4241 997 -4195 1009
rect -4241 121 -4235 997
rect -4201 121 -4195 997
rect -4241 109 -4195 121
rect -4093 997 -4047 1009
rect -4093 121 -4087 997
rect -4053 121 -4047 997
rect -4093 109 -4047 121
rect -3945 997 -3899 1009
rect -3945 121 -3939 997
rect -3905 121 -3899 997
rect -3945 109 -3899 121
rect -3797 997 -3751 1009
rect -3797 121 -3791 997
rect -3757 121 -3751 997
rect -3797 109 -3751 121
rect -3649 997 -3603 1009
rect -3649 121 -3643 997
rect -3609 121 -3603 997
rect -3649 109 -3603 121
rect -3501 997 -3455 1009
rect -3501 121 -3495 997
rect -3461 121 -3455 997
rect -3501 109 -3455 121
rect -3353 997 -3307 1009
rect -3353 121 -3347 997
rect -3313 121 -3307 997
rect -3353 109 -3307 121
rect -3205 997 -3159 1009
rect -3205 121 -3199 997
rect -3165 121 -3159 997
rect -3205 109 -3159 121
rect -3057 997 -3011 1009
rect -3057 121 -3051 997
rect -3017 121 -3011 997
rect -3057 109 -3011 121
rect -2909 997 -2863 1009
rect -2909 121 -2903 997
rect -2869 121 -2863 997
rect -2909 109 -2863 121
rect -2761 997 -2715 1009
rect -2761 121 -2755 997
rect -2721 121 -2715 997
rect -2761 109 -2715 121
rect -2613 997 -2567 1009
rect -2613 121 -2607 997
rect -2573 121 -2567 997
rect -2613 109 -2567 121
rect -2465 997 -2419 1009
rect -2465 121 -2459 997
rect -2425 121 -2419 997
rect -2465 109 -2419 121
rect -2317 997 -2271 1009
rect -2317 121 -2311 997
rect -2277 121 -2271 997
rect -2317 109 -2271 121
rect -2169 997 -2123 1009
rect -2169 121 -2163 997
rect -2129 121 -2123 997
rect -2169 109 -2123 121
rect -2021 997 -1975 1009
rect -2021 121 -2015 997
rect -1981 121 -1975 997
rect -2021 109 -1975 121
rect -1873 997 -1827 1009
rect -1873 121 -1867 997
rect -1833 121 -1827 997
rect -1873 109 -1827 121
rect -1725 997 -1679 1009
rect -1725 121 -1719 997
rect -1685 121 -1679 997
rect -1725 109 -1679 121
rect -1577 997 -1531 1009
rect -1577 121 -1571 997
rect -1537 121 -1531 997
rect -1577 109 -1531 121
rect -1429 997 -1383 1009
rect -1429 121 -1423 997
rect -1389 121 -1383 997
rect -1429 109 -1383 121
rect -1281 997 -1235 1009
rect -1281 121 -1275 997
rect -1241 121 -1235 997
rect -1281 109 -1235 121
rect -1133 997 -1087 1009
rect -1133 121 -1127 997
rect -1093 121 -1087 997
rect -1133 109 -1087 121
rect -985 997 -939 1009
rect -985 121 -979 997
rect -945 121 -939 997
rect -985 109 -939 121
rect -837 997 -791 1009
rect -837 121 -831 997
rect -797 121 -791 997
rect -837 109 -791 121
rect -689 997 -643 1009
rect -689 121 -683 997
rect -649 121 -643 997
rect -689 109 -643 121
rect -541 997 -495 1009
rect -541 121 -535 997
rect -501 121 -495 997
rect -541 109 -495 121
rect -393 997 -347 1009
rect -393 121 -387 997
rect -353 121 -347 997
rect -393 109 -347 121
rect -245 997 -199 1009
rect -245 121 -239 997
rect -205 121 -199 997
rect -245 109 -199 121
rect -97 997 -51 1009
rect -97 121 -91 997
rect -57 121 -51 997
rect -97 109 -51 121
rect 51 997 97 1009
rect 51 121 57 997
rect 91 121 97 997
rect 51 109 97 121
rect 199 997 245 1009
rect 199 121 205 997
rect 239 121 245 997
rect 199 109 245 121
rect 347 997 393 1009
rect 347 121 353 997
rect 387 121 393 997
rect 347 109 393 121
rect 495 997 541 1009
rect 495 121 501 997
rect 535 121 541 997
rect 495 109 541 121
rect 643 997 689 1009
rect 643 121 649 997
rect 683 121 689 997
rect 643 109 689 121
rect 791 997 837 1009
rect 791 121 797 997
rect 831 121 837 997
rect 791 109 837 121
rect 939 997 985 1009
rect 939 121 945 997
rect 979 121 985 997
rect 939 109 985 121
rect 1087 997 1133 1009
rect 1087 121 1093 997
rect 1127 121 1133 997
rect 1087 109 1133 121
rect 1235 997 1281 1009
rect 1235 121 1241 997
rect 1275 121 1281 997
rect 1235 109 1281 121
rect 1383 997 1429 1009
rect 1383 121 1389 997
rect 1423 121 1429 997
rect 1383 109 1429 121
rect 1531 997 1577 1009
rect 1531 121 1537 997
rect 1571 121 1577 997
rect 1531 109 1577 121
rect 1679 997 1725 1009
rect 1679 121 1685 997
rect 1719 121 1725 997
rect 1679 109 1725 121
rect 1827 997 1873 1009
rect 1827 121 1833 997
rect 1867 121 1873 997
rect 1827 109 1873 121
rect 1975 997 2021 1009
rect 1975 121 1981 997
rect 2015 121 2021 997
rect 1975 109 2021 121
rect 2123 997 2169 1009
rect 2123 121 2129 997
rect 2163 121 2169 997
rect 2123 109 2169 121
rect 2271 997 2317 1009
rect 2271 121 2277 997
rect 2311 121 2317 997
rect 2271 109 2317 121
rect 2419 997 2465 1009
rect 2419 121 2425 997
rect 2459 121 2465 997
rect 2419 109 2465 121
rect 2567 997 2613 1009
rect 2567 121 2573 997
rect 2607 121 2613 997
rect 2567 109 2613 121
rect 2715 997 2761 1009
rect 2715 121 2721 997
rect 2755 121 2761 997
rect 2715 109 2761 121
rect 2863 997 2909 1009
rect 2863 121 2869 997
rect 2903 121 2909 997
rect 2863 109 2909 121
rect 3011 997 3057 1009
rect 3011 121 3017 997
rect 3051 121 3057 997
rect 3011 109 3057 121
rect 3159 997 3205 1009
rect 3159 121 3165 997
rect 3199 121 3205 997
rect 3159 109 3205 121
rect 3307 997 3353 1009
rect 3307 121 3313 997
rect 3347 121 3353 997
rect 3307 109 3353 121
rect 3455 997 3501 1009
rect 3455 121 3461 997
rect 3495 121 3501 997
rect 3455 109 3501 121
rect 3603 997 3649 1009
rect 3603 121 3609 997
rect 3643 121 3649 997
rect 3603 109 3649 121
rect 3751 997 3797 1009
rect 3751 121 3757 997
rect 3791 121 3797 997
rect 3751 109 3797 121
rect 3899 997 3945 1009
rect 3899 121 3905 997
rect 3939 121 3945 997
rect 3899 109 3945 121
rect 4047 997 4093 1009
rect 4047 121 4053 997
rect 4087 121 4093 997
rect 4047 109 4093 121
rect 4195 997 4241 1009
rect 4195 121 4201 997
rect 4235 121 4241 997
rect 4195 109 4241 121
rect 4343 997 4389 1009
rect 4343 121 4349 997
rect 4383 121 4389 997
rect 4343 109 4389 121
rect 4491 997 4537 1009
rect 4491 121 4497 997
rect 4531 121 4537 997
rect 4491 109 4537 121
rect 4639 997 4685 1009
rect 4639 121 4645 997
rect 4679 121 4685 997
rect 4639 109 4685 121
rect 4787 997 4833 1009
rect 4787 121 4793 997
rect 4827 121 4833 997
rect 4787 109 4833 121
rect 4935 997 4981 1009
rect 4935 121 4941 997
rect 4975 121 4981 997
rect 4935 109 4981 121
rect 5083 997 5129 1009
rect 5083 121 5089 997
rect 5123 121 5129 997
rect 5083 109 5129 121
rect 5231 997 5277 1009
rect 5231 121 5237 997
rect 5271 121 5277 997
rect 5231 109 5277 121
rect 5379 997 5425 1009
rect 5379 121 5385 997
rect 5419 121 5425 997
rect 5379 109 5425 121
rect 5527 997 5573 1009
rect 5527 121 5533 997
rect 5567 121 5573 997
rect 5527 109 5573 121
rect -5517 71 -5435 77
rect -5517 37 -5505 71
rect -5447 37 -5435 71
rect -5517 31 -5435 37
rect -5369 71 -5287 77
rect -5369 37 -5357 71
rect -5299 37 -5287 71
rect -5369 31 -5287 37
rect -5221 71 -5139 77
rect -5221 37 -5209 71
rect -5151 37 -5139 71
rect -5221 31 -5139 37
rect -5073 71 -4991 77
rect -5073 37 -5061 71
rect -5003 37 -4991 71
rect -5073 31 -4991 37
rect -4925 71 -4843 77
rect -4925 37 -4913 71
rect -4855 37 -4843 71
rect -4925 31 -4843 37
rect -4777 71 -4695 77
rect -4777 37 -4765 71
rect -4707 37 -4695 71
rect -4777 31 -4695 37
rect -4629 71 -4547 77
rect -4629 37 -4617 71
rect -4559 37 -4547 71
rect -4629 31 -4547 37
rect -4481 71 -4399 77
rect -4481 37 -4469 71
rect -4411 37 -4399 71
rect -4481 31 -4399 37
rect -4333 71 -4251 77
rect -4333 37 -4321 71
rect -4263 37 -4251 71
rect -4333 31 -4251 37
rect -4185 71 -4103 77
rect -4185 37 -4173 71
rect -4115 37 -4103 71
rect -4185 31 -4103 37
rect -4037 71 -3955 77
rect -4037 37 -4025 71
rect -3967 37 -3955 71
rect -4037 31 -3955 37
rect -3889 71 -3807 77
rect -3889 37 -3877 71
rect -3819 37 -3807 71
rect -3889 31 -3807 37
rect -3741 71 -3659 77
rect -3741 37 -3729 71
rect -3671 37 -3659 71
rect -3741 31 -3659 37
rect -3593 71 -3511 77
rect -3593 37 -3581 71
rect -3523 37 -3511 71
rect -3593 31 -3511 37
rect -3445 71 -3363 77
rect -3445 37 -3433 71
rect -3375 37 -3363 71
rect -3445 31 -3363 37
rect -3297 71 -3215 77
rect -3297 37 -3285 71
rect -3227 37 -3215 71
rect -3297 31 -3215 37
rect -3149 71 -3067 77
rect -3149 37 -3137 71
rect -3079 37 -3067 71
rect -3149 31 -3067 37
rect -3001 71 -2919 77
rect -3001 37 -2989 71
rect -2931 37 -2919 71
rect -3001 31 -2919 37
rect -2853 71 -2771 77
rect -2853 37 -2841 71
rect -2783 37 -2771 71
rect -2853 31 -2771 37
rect -2705 71 -2623 77
rect -2705 37 -2693 71
rect -2635 37 -2623 71
rect -2705 31 -2623 37
rect -2557 71 -2475 77
rect -2557 37 -2545 71
rect -2487 37 -2475 71
rect -2557 31 -2475 37
rect -2409 71 -2327 77
rect -2409 37 -2397 71
rect -2339 37 -2327 71
rect -2409 31 -2327 37
rect -2261 71 -2179 77
rect -2261 37 -2249 71
rect -2191 37 -2179 71
rect -2261 31 -2179 37
rect -2113 71 -2031 77
rect -2113 37 -2101 71
rect -2043 37 -2031 71
rect -2113 31 -2031 37
rect -1965 71 -1883 77
rect -1965 37 -1953 71
rect -1895 37 -1883 71
rect -1965 31 -1883 37
rect -1817 71 -1735 77
rect -1817 37 -1805 71
rect -1747 37 -1735 71
rect -1817 31 -1735 37
rect -1669 71 -1587 77
rect -1669 37 -1657 71
rect -1599 37 -1587 71
rect -1669 31 -1587 37
rect -1521 71 -1439 77
rect -1521 37 -1509 71
rect -1451 37 -1439 71
rect -1521 31 -1439 37
rect -1373 71 -1291 77
rect -1373 37 -1361 71
rect -1303 37 -1291 71
rect -1373 31 -1291 37
rect -1225 71 -1143 77
rect -1225 37 -1213 71
rect -1155 37 -1143 71
rect -1225 31 -1143 37
rect -1077 71 -995 77
rect -1077 37 -1065 71
rect -1007 37 -995 71
rect -1077 31 -995 37
rect -929 71 -847 77
rect -929 37 -917 71
rect -859 37 -847 71
rect -929 31 -847 37
rect -781 71 -699 77
rect -781 37 -769 71
rect -711 37 -699 71
rect -781 31 -699 37
rect -633 71 -551 77
rect -633 37 -621 71
rect -563 37 -551 71
rect -633 31 -551 37
rect -485 71 -403 77
rect -485 37 -473 71
rect -415 37 -403 71
rect -485 31 -403 37
rect -337 71 -255 77
rect -337 37 -325 71
rect -267 37 -255 71
rect -337 31 -255 37
rect -189 71 -107 77
rect -189 37 -177 71
rect -119 37 -107 71
rect -189 31 -107 37
rect -41 71 41 77
rect -41 37 -29 71
rect 29 37 41 71
rect -41 31 41 37
rect 107 71 189 77
rect 107 37 119 71
rect 177 37 189 71
rect 107 31 189 37
rect 255 71 337 77
rect 255 37 267 71
rect 325 37 337 71
rect 255 31 337 37
rect 403 71 485 77
rect 403 37 415 71
rect 473 37 485 71
rect 403 31 485 37
rect 551 71 633 77
rect 551 37 563 71
rect 621 37 633 71
rect 551 31 633 37
rect 699 71 781 77
rect 699 37 711 71
rect 769 37 781 71
rect 699 31 781 37
rect 847 71 929 77
rect 847 37 859 71
rect 917 37 929 71
rect 847 31 929 37
rect 995 71 1077 77
rect 995 37 1007 71
rect 1065 37 1077 71
rect 995 31 1077 37
rect 1143 71 1225 77
rect 1143 37 1155 71
rect 1213 37 1225 71
rect 1143 31 1225 37
rect 1291 71 1373 77
rect 1291 37 1303 71
rect 1361 37 1373 71
rect 1291 31 1373 37
rect 1439 71 1521 77
rect 1439 37 1451 71
rect 1509 37 1521 71
rect 1439 31 1521 37
rect 1587 71 1669 77
rect 1587 37 1599 71
rect 1657 37 1669 71
rect 1587 31 1669 37
rect 1735 71 1817 77
rect 1735 37 1747 71
rect 1805 37 1817 71
rect 1735 31 1817 37
rect 1883 71 1965 77
rect 1883 37 1895 71
rect 1953 37 1965 71
rect 1883 31 1965 37
rect 2031 71 2113 77
rect 2031 37 2043 71
rect 2101 37 2113 71
rect 2031 31 2113 37
rect 2179 71 2261 77
rect 2179 37 2191 71
rect 2249 37 2261 71
rect 2179 31 2261 37
rect 2327 71 2409 77
rect 2327 37 2339 71
rect 2397 37 2409 71
rect 2327 31 2409 37
rect 2475 71 2557 77
rect 2475 37 2487 71
rect 2545 37 2557 71
rect 2475 31 2557 37
rect 2623 71 2705 77
rect 2623 37 2635 71
rect 2693 37 2705 71
rect 2623 31 2705 37
rect 2771 71 2853 77
rect 2771 37 2783 71
rect 2841 37 2853 71
rect 2771 31 2853 37
rect 2919 71 3001 77
rect 2919 37 2931 71
rect 2989 37 3001 71
rect 2919 31 3001 37
rect 3067 71 3149 77
rect 3067 37 3079 71
rect 3137 37 3149 71
rect 3067 31 3149 37
rect 3215 71 3297 77
rect 3215 37 3227 71
rect 3285 37 3297 71
rect 3215 31 3297 37
rect 3363 71 3445 77
rect 3363 37 3375 71
rect 3433 37 3445 71
rect 3363 31 3445 37
rect 3511 71 3593 77
rect 3511 37 3523 71
rect 3581 37 3593 71
rect 3511 31 3593 37
rect 3659 71 3741 77
rect 3659 37 3671 71
rect 3729 37 3741 71
rect 3659 31 3741 37
rect 3807 71 3889 77
rect 3807 37 3819 71
rect 3877 37 3889 71
rect 3807 31 3889 37
rect 3955 71 4037 77
rect 3955 37 3967 71
rect 4025 37 4037 71
rect 3955 31 4037 37
rect 4103 71 4185 77
rect 4103 37 4115 71
rect 4173 37 4185 71
rect 4103 31 4185 37
rect 4251 71 4333 77
rect 4251 37 4263 71
rect 4321 37 4333 71
rect 4251 31 4333 37
rect 4399 71 4481 77
rect 4399 37 4411 71
rect 4469 37 4481 71
rect 4399 31 4481 37
rect 4547 71 4629 77
rect 4547 37 4559 71
rect 4617 37 4629 71
rect 4547 31 4629 37
rect 4695 71 4777 77
rect 4695 37 4707 71
rect 4765 37 4777 71
rect 4695 31 4777 37
rect 4843 71 4925 77
rect 4843 37 4855 71
rect 4913 37 4925 71
rect 4843 31 4925 37
rect 4991 71 5073 77
rect 4991 37 5003 71
rect 5061 37 5073 71
rect 4991 31 5073 37
rect 5139 71 5221 77
rect 5139 37 5151 71
rect 5209 37 5221 71
rect 5139 31 5221 37
rect 5287 71 5369 77
rect 5287 37 5299 71
rect 5357 37 5369 71
rect 5287 31 5369 37
rect 5435 71 5517 77
rect 5435 37 5447 71
rect 5505 37 5517 71
rect 5435 31 5517 37
rect -5517 -37 -5435 -31
rect -5517 -71 -5505 -37
rect -5447 -71 -5435 -37
rect -5517 -77 -5435 -71
rect -5369 -37 -5287 -31
rect -5369 -71 -5357 -37
rect -5299 -71 -5287 -37
rect -5369 -77 -5287 -71
rect -5221 -37 -5139 -31
rect -5221 -71 -5209 -37
rect -5151 -71 -5139 -37
rect -5221 -77 -5139 -71
rect -5073 -37 -4991 -31
rect -5073 -71 -5061 -37
rect -5003 -71 -4991 -37
rect -5073 -77 -4991 -71
rect -4925 -37 -4843 -31
rect -4925 -71 -4913 -37
rect -4855 -71 -4843 -37
rect -4925 -77 -4843 -71
rect -4777 -37 -4695 -31
rect -4777 -71 -4765 -37
rect -4707 -71 -4695 -37
rect -4777 -77 -4695 -71
rect -4629 -37 -4547 -31
rect -4629 -71 -4617 -37
rect -4559 -71 -4547 -37
rect -4629 -77 -4547 -71
rect -4481 -37 -4399 -31
rect -4481 -71 -4469 -37
rect -4411 -71 -4399 -37
rect -4481 -77 -4399 -71
rect -4333 -37 -4251 -31
rect -4333 -71 -4321 -37
rect -4263 -71 -4251 -37
rect -4333 -77 -4251 -71
rect -4185 -37 -4103 -31
rect -4185 -71 -4173 -37
rect -4115 -71 -4103 -37
rect -4185 -77 -4103 -71
rect -4037 -37 -3955 -31
rect -4037 -71 -4025 -37
rect -3967 -71 -3955 -37
rect -4037 -77 -3955 -71
rect -3889 -37 -3807 -31
rect -3889 -71 -3877 -37
rect -3819 -71 -3807 -37
rect -3889 -77 -3807 -71
rect -3741 -37 -3659 -31
rect -3741 -71 -3729 -37
rect -3671 -71 -3659 -37
rect -3741 -77 -3659 -71
rect -3593 -37 -3511 -31
rect -3593 -71 -3581 -37
rect -3523 -71 -3511 -37
rect -3593 -77 -3511 -71
rect -3445 -37 -3363 -31
rect -3445 -71 -3433 -37
rect -3375 -71 -3363 -37
rect -3445 -77 -3363 -71
rect -3297 -37 -3215 -31
rect -3297 -71 -3285 -37
rect -3227 -71 -3215 -37
rect -3297 -77 -3215 -71
rect -3149 -37 -3067 -31
rect -3149 -71 -3137 -37
rect -3079 -71 -3067 -37
rect -3149 -77 -3067 -71
rect -3001 -37 -2919 -31
rect -3001 -71 -2989 -37
rect -2931 -71 -2919 -37
rect -3001 -77 -2919 -71
rect -2853 -37 -2771 -31
rect -2853 -71 -2841 -37
rect -2783 -71 -2771 -37
rect -2853 -77 -2771 -71
rect -2705 -37 -2623 -31
rect -2705 -71 -2693 -37
rect -2635 -71 -2623 -37
rect -2705 -77 -2623 -71
rect -2557 -37 -2475 -31
rect -2557 -71 -2545 -37
rect -2487 -71 -2475 -37
rect -2557 -77 -2475 -71
rect -2409 -37 -2327 -31
rect -2409 -71 -2397 -37
rect -2339 -71 -2327 -37
rect -2409 -77 -2327 -71
rect -2261 -37 -2179 -31
rect -2261 -71 -2249 -37
rect -2191 -71 -2179 -37
rect -2261 -77 -2179 -71
rect -2113 -37 -2031 -31
rect -2113 -71 -2101 -37
rect -2043 -71 -2031 -37
rect -2113 -77 -2031 -71
rect -1965 -37 -1883 -31
rect -1965 -71 -1953 -37
rect -1895 -71 -1883 -37
rect -1965 -77 -1883 -71
rect -1817 -37 -1735 -31
rect -1817 -71 -1805 -37
rect -1747 -71 -1735 -37
rect -1817 -77 -1735 -71
rect -1669 -37 -1587 -31
rect -1669 -71 -1657 -37
rect -1599 -71 -1587 -37
rect -1669 -77 -1587 -71
rect -1521 -37 -1439 -31
rect -1521 -71 -1509 -37
rect -1451 -71 -1439 -37
rect -1521 -77 -1439 -71
rect -1373 -37 -1291 -31
rect -1373 -71 -1361 -37
rect -1303 -71 -1291 -37
rect -1373 -77 -1291 -71
rect -1225 -37 -1143 -31
rect -1225 -71 -1213 -37
rect -1155 -71 -1143 -37
rect -1225 -77 -1143 -71
rect -1077 -37 -995 -31
rect -1077 -71 -1065 -37
rect -1007 -71 -995 -37
rect -1077 -77 -995 -71
rect -929 -37 -847 -31
rect -929 -71 -917 -37
rect -859 -71 -847 -37
rect -929 -77 -847 -71
rect -781 -37 -699 -31
rect -781 -71 -769 -37
rect -711 -71 -699 -37
rect -781 -77 -699 -71
rect -633 -37 -551 -31
rect -633 -71 -621 -37
rect -563 -71 -551 -37
rect -633 -77 -551 -71
rect -485 -37 -403 -31
rect -485 -71 -473 -37
rect -415 -71 -403 -37
rect -485 -77 -403 -71
rect -337 -37 -255 -31
rect -337 -71 -325 -37
rect -267 -71 -255 -37
rect -337 -77 -255 -71
rect -189 -37 -107 -31
rect -189 -71 -177 -37
rect -119 -71 -107 -37
rect -189 -77 -107 -71
rect -41 -37 41 -31
rect -41 -71 -29 -37
rect 29 -71 41 -37
rect -41 -77 41 -71
rect 107 -37 189 -31
rect 107 -71 119 -37
rect 177 -71 189 -37
rect 107 -77 189 -71
rect 255 -37 337 -31
rect 255 -71 267 -37
rect 325 -71 337 -37
rect 255 -77 337 -71
rect 403 -37 485 -31
rect 403 -71 415 -37
rect 473 -71 485 -37
rect 403 -77 485 -71
rect 551 -37 633 -31
rect 551 -71 563 -37
rect 621 -71 633 -37
rect 551 -77 633 -71
rect 699 -37 781 -31
rect 699 -71 711 -37
rect 769 -71 781 -37
rect 699 -77 781 -71
rect 847 -37 929 -31
rect 847 -71 859 -37
rect 917 -71 929 -37
rect 847 -77 929 -71
rect 995 -37 1077 -31
rect 995 -71 1007 -37
rect 1065 -71 1077 -37
rect 995 -77 1077 -71
rect 1143 -37 1225 -31
rect 1143 -71 1155 -37
rect 1213 -71 1225 -37
rect 1143 -77 1225 -71
rect 1291 -37 1373 -31
rect 1291 -71 1303 -37
rect 1361 -71 1373 -37
rect 1291 -77 1373 -71
rect 1439 -37 1521 -31
rect 1439 -71 1451 -37
rect 1509 -71 1521 -37
rect 1439 -77 1521 -71
rect 1587 -37 1669 -31
rect 1587 -71 1599 -37
rect 1657 -71 1669 -37
rect 1587 -77 1669 -71
rect 1735 -37 1817 -31
rect 1735 -71 1747 -37
rect 1805 -71 1817 -37
rect 1735 -77 1817 -71
rect 1883 -37 1965 -31
rect 1883 -71 1895 -37
rect 1953 -71 1965 -37
rect 1883 -77 1965 -71
rect 2031 -37 2113 -31
rect 2031 -71 2043 -37
rect 2101 -71 2113 -37
rect 2031 -77 2113 -71
rect 2179 -37 2261 -31
rect 2179 -71 2191 -37
rect 2249 -71 2261 -37
rect 2179 -77 2261 -71
rect 2327 -37 2409 -31
rect 2327 -71 2339 -37
rect 2397 -71 2409 -37
rect 2327 -77 2409 -71
rect 2475 -37 2557 -31
rect 2475 -71 2487 -37
rect 2545 -71 2557 -37
rect 2475 -77 2557 -71
rect 2623 -37 2705 -31
rect 2623 -71 2635 -37
rect 2693 -71 2705 -37
rect 2623 -77 2705 -71
rect 2771 -37 2853 -31
rect 2771 -71 2783 -37
rect 2841 -71 2853 -37
rect 2771 -77 2853 -71
rect 2919 -37 3001 -31
rect 2919 -71 2931 -37
rect 2989 -71 3001 -37
rect 2919 -77 3001 -71
rect 3067 -37 3149 -31
rect 3067 -71 3079 -37
rect 3137 -71 3149 -37
rect 3067 -77 3149 -71
rect 3215 -37 3297 -31
rect 3215 -71 3227 -37
rect 3285 -71 3297 -37
rect 3215 -77 3297 -71
rect 3363 -37 3445 -31
rect 3363 -71 3375 -37
rect 3433 -71 3445 -37
rect 3363 -77 3445 -71
rect 3511 -37 3593 -31
rect 3511 -71 3523 -37
rect 3581 -71 3593 -37
rect 3511 -77 3593 -71
rect 3659 -37 3741 -31
rect 3659 -71 3671 -37
rect 3729 -71 3741 -37
rect 3659 -77 3741 -71
rect 3807 -37 3889 -31
rect 3807 -71 3819 -37
rect 3877 -71 3889 -37
rect 3807 -77 3889 -71
rect 3955 -37 4037 -31
rect 3955 -71 3967 -37
rect 4025 -71 4037 -37
rect 3955 -77 4037 -71
rect 4103 -37 4185 -31
rect 4103 -71 4115 -37
rect 4173 -71 4185 -37
rect 4103 -77 4185 -71
rect 4251 -37 4333 -31
rect 4251 -71 4263 -37
rect 4321 -71 4333 -37
rect 4251 -77 4333 -71
rect 4399 -37 4481 -31
rect 4399 -71 4411 -37
rect 4469 -71 4481 -37
rect 4399 -77 4481 -71
rect 4547 -37 4629 -31
rect 4547 -71 4559 -37
rect 4617 -71 4629 -37
rect 4547 -77 4629 -71
rect 4695 -37 4777 -31
rect 4695 -71 4707 -37
rect 4765 -71 4777 -37
rect 4695 -77 4777 -71
rect 4843 -37 4925 -31
rect 4843 -71 4855 -37
rect 4913 -71 4925 -37
rect 4843 -77 4925 -71
rect 4991 -37 5073 -31
rect 4991 -71 5003 -37
rect 5061 -71 5073 -37
rect 4991 -77 5073 -71
rect 5139 -37 5221 -31
rect 5139 -71 5151 -37
rect 5209 -71 5221 -37
rect 5139 -77 5221 -71
rect 5287 -37 5369 -31
rect 5287 -71 5299 -37
rect 5357 -71 5369 -37
rect 5287 -77 5369 -71
rect 5435 -37 5517 -31
rect 5435 -71 5447 -37
rect 5505 -71 5517 -37
rect 5435 -77 5517 -71
rect -5573 -121 -5527 -109
rect -5573 -997 -5567 -121
rect -5533 -997 -5527 -121
rect -5573 -1009 -5527 -997
rect -5425 -121 -5379 -109
rect -5425 -997 -5419 -121
rect -5385 -997 -5379 -121
rect -5425 -1009 -5379 -997
rect -5277 -121 -5231 -109
rect -5277 -997 -5271 -121
rect -5237 -997 -5231 -121
rect -5277 -1009 -5231 -997
rect -5129 -121 -5083 -109
rect -5129 -997 -5123 -121
rect -5089 -997 -5083 -121
rect -5129 -1009 -5083 -997
rect -4981 -121 -4935 -109
rect -4981 -997 -4975 -121
rect -4941 -997 -4935 -121
rect -4981 -1009 -4935 -997
rect -4833 -121 -4787 -109
rect -4833 -997 -4827 -121
rect -4793 -997 -4787 -121
rect -4833 -1009 -4787 -997
rect -4685 -121 -4639 -109
rect -4685 -997 -4679 -121
rect -4645 -997 -4639 -121
rect -4685 -1009 -4639 -997
rect -4537 -121 -4491 -109
rect -4537 -997 -4531 -121
rect -4497 -997 -4491 -121
rect -4537 -1009 -4491 -997
rect -4389 -121 -4343 -109
rect -4389 -997 -4383 -121
rect -4349 -997 -4343 -121
rect -4389 -1009 -4343 -997
rect -4241 -121 -4195 -109
rect -4241 -997 -4235 -121
rect -4201 -997 -4195 -121
rect -4241 -1009 -4195 -997
rect -4093 -121 -4047 -109
rect -4093 -997 -4087 -121
rect -4053 -997 -4047 -121
rect -4093 -1009 -4047 -997
rect -3945 -121 -3899 -109
rect -3945 -997 -3939 -121
rect -3905 -997 -3899 -121
rect -3945 -1009 -3899 -997
rect -3797 -121 -3751 -109
rect -3797 -997 -3791 -121
rect -3757 -997 -3751 -121
rect -3797 -1009 -3751 -997
rect -3649 -121 -3603 -109
rect -3649 -997 -3643 -121
rect -3609 -997 -3603 -121
rect -3649 -1009 -3603 -997
rect -3501 -121 -3455 -109
rect -3501 -997 -3495 -121
rect -3461 -997 -3455 -121
rect -3501 -1009 -3455 -997
rect -3353 -121 -3307 -109
rect -3353 -997 -3347 -121
rect -3313 -997 -3307 -121
rect -3353 -1009 -3307 -997
rect -3205 -121 -3159 -109
rect -3205 -997 -3199 -121
rect -3165 -997 -3159 -121
rect -3205 -1009 -3159 -997
rect -3057 -121 -3011 -109
rect -3057 -997 -3051 -121
rect -3017 -997 -3011 -121
rect -3057 -1009 -3011 -997
rect -2909 -121 -2863 -109
rect -2909 -997 -2903 -121
rect -2869 -997 -2863 -121
rect -2909 -1009 -2863 -997
rect -2761 -121 -2715 -109
rect -2761 -997 -2755 -121
rect -2721 -997 -2715 -121
rect -2761 -1009 -2715 -997
rect -2613 -121 -2567 -109
rect -2613 -997 -2607 -121
rect -2573 -997 -2567 -121
rect -2613 -1009 -2567 -997
rect -2465 -121 -2419 -109
rect -2465 -997 -2459 -121
rect -2425 -997 -2419 -121
rect -2465 -1009 -2419 -997
rect -2317 -121 -2271 -109
rect -2317 -997 -2311 -121
rect -2277 -997 -2271 -121
rect -2317 -1009 -2271 -997
rect -2169 -121 -2123 -109
rect -2169 -997 -2163 -121
rect -2129 -997 -2123 -121
rect -2169 -1009 -2123 -997
rect -2021 -121 -1975 -109
rect -2021 -997 -2015 -121
rect -1981 -997 -1975 -121
rect -2021 -1009 -1975 -997
rect -1873 -121 -1827 -109
rect -1873 -997 -1867 -121
rect -1833 -997 -1827 -121
rect -1873 -1009 -1827 -997
rect -1725 -121 -1679 -109
rect -1725 -997 -1719 -121
rect -1685 -997 -1679 -121
rect -1725 -1009 -1679 -997
rect -1577 -121 -1531 -109
rect -1577 -997 -1571 -121
rect -1537 -997 -1531 -121
rect -1577 -1009 -1531 -997
rect -1429 -121 -1383 -109
rect -1429 -997 -1423 -121
rect -1389 -997 -1383 -121
rect -1429 -1009 -1383 -997
rect -1281 -121 -1235 -109
rect -1281 -997 -1275 -121
rect -1241 -997 -1235 -121
rect -1281 -1009 -1235 -997
rect -1133 -121 -1087 -109
rect -1133 -997 -1127 -121
rect -1093 -997 -1087 -121
rect -1133 -1009 -1087 -997
rect -985 -121 -939 -109
rect -985 -997 -979 -121
rect -945 -997 -939 -121
rect -985 -1009 -939 -997
rect -837 -121 -791 -109
rect -837 -997 -831 -121
rect -797 -997 -791 -121
rect -837 -1009 -791 -997
rect -689 -121 -643 -109
rect -689 -997 -683 -121
rect -649 -997 -643 -121
rect -689 -1009 -643 -997
rect -541 -121 -495 -109
rect -541 -997 -535 -121
rect -501 -997 -495 -121
rect -541 -1009 -495 -997
rect -393 -121 -347 -109
rect -393 -997 -387 -121
rect -353 -997 -347 -121
rect -393 -1009 -347 -997
rect -245 -121 -199 -109
rect -245 -997 -239 -121
rect -205 -997 -199 -121
rect -245 -1009 -199 -997
rect -97 -121 -51 -109
rect -97 -997 -91 -121
rect -57 -997 -51 -121
rect -97 -1009 -51 -997
rect 51 -121 97 -109
rect 51 -997 57 -121
rect 91 -997 97 -121
rect 51 -1009 97 -997
rect 199 -121 245 -109
rect 199 -997 205 -121
rect 239 -997 245 -121
rect 199 -1009 245 -997
rect 347 -121 393 -109
rect 347 -997 353 -121
rect 387 -997 393 -121
rect 347 -1009 393 -997
rect 495 -121 541 -109
rect 495 -997 501 -121
rect 535 -997 541 -121
rect 495 -1009 541 -997
rect 643 -121 689 -109
rect 643 -997 649 -121
rect 683 -997 689 -121
rect 643 -1009 689 -997
rect 791 -121 837 -109
rect 791 -997 797 -121
rect 831 -997 837 -121
rect 791 -1009 837 -997
rect 939 -121 985 -109
rect 939 -997 945 -121
rect 979 -997 985 -121
rect 939 -1009 985 -997
rect 1087 -121 1133 -109
rect 1087 -997 1093 -121
rect 1127 -997 1133 -121
rect 1087 -1009 1133 -997
rect 1235 -121 1281 -109
rect 1235 -997 1241 -121
rect 1275 -997 1281 -121
rect 1235 -1009 1281 -997
rect 1383 -121 1429 -109
rect 1383 -997 1389 -121
rect 1423 -997 1429 -121
rect 1383 -1009 1429 -997
rect 1531 -121 1577 -109
rect 1531 -997 1537 -121
rect 1571 -997 1577 -121
rect 1531 -1009 1577 -997
rect 1679 -121 1725 -109
rect 1679 -997 1685 -121
rect 1719 -997 1725 -121
rect 1679 -1009 1725 -997
rect 1827 -121 1873 -109
rect 1827 -997 1833 -121
rect 1867 -997 1873 -121
rect 1827 -1009 1873 -997
rect 1975 -121 2021 -109
rect 1975 -997 1981 -121
rect 2015 -997 2021 -121
rect 1975 -1009 2021 -997
rect 2123 -121 2169 -109
rect 2123 -997 2129 -121
rect 2163 -997 2169 -121
rect 2123 -1009 2169 -997
rect 2271 -121 2317 -109
rect 2271 -997 2277 -121
rect 2311 -997 2317 -121
rect 2271 -1009 2317 -997
rect 2419 -121 2465 -109
rect 2419 -997 2425 -121
rect 2459 -997 2465 -121
rect 2419 -1009 2465 -997
rect 2567 -121 2613 -109
rect 2567 -997 2573 -121
rect 2607 -997 2613 -121
rect 2567 -1009 2613 -997
rect 2715 -121 2761 -109
rect 2715 -997 2721 -121
rect 2755 -997 2761 -121
rect 2715 -1009 2761 -997
rect 2863 -121 2909 -109
rect 2863 -997 2869 -121
rect 2903 -997 2909 -121
rect 2863 -1009 2909 -997
rect 3011 -121 3057 -109
rect 3011 -997 3017 -121
rect 3051 -997 3057 -121
rect 3011 -1009 3057 -997
rect 3159 -121 3205 -109
rect 3159 -997 3165 -121
rect 3199 -997 3205 -121
rect 3159 -1009 3205 -997
rect 3307 -121 3353 -109
rect 3307 -997 3313 -121
rect 3347 -997 3353 -121
rect 3307 -1009 3353 -997
rect 3455 -121 3501 -109
rect 3455 -997 3461 -121
rect 3495 -997 3501 -121
rect 3455 -1009 3501 -997
rect 3603 -121 3649 -109
rect 3603 -997 3609 -121
rect 3643 -997 3649 -121
rect 3603 -1009 3649 -997
rect 3751 -121 3797 -109
rect 3751 -997 3757 -121
rect 3791 -997 3797 -121
rect 3751 -1009 3797 -997
rect 3899 -121 3945 -109
rect 3899 -997 3905 -121
rect 3939 -997 3945 -121
rect 3899 -1009 3945 -997
rect 4047 -121 4093 -109
rect 4047 -997 4053 -121
rect 4087 -997 4093 -121
rect 4047 -1009 4093 -997
rect 4195 -121 4241 -109
rect 4195 -997 4201 -121
rect 4235 -997 4241 -121
rect 4195 -1009 4241 -997
rect 4343 -121 4389 -109
rect 4343 -997 4349 -121
rect 4383 -997 4389 -121
rect 4343 -1009 4389 -997
rect 4491 -121 4537 -109
rect 4491 -997 4497 -121
rect 4531 -997 4537 -121
rect 4491 -1009 4537 -997
rect 4639 -121 4685 -109
rect 4639 -997 4645 -121
rect 4679 -997 4685 -121
rect 4639 -1009 4685 -997
rect 4787 -121 4833 -109
rect 4787 -997 4793 -121
rect 4827 -997 4833 -121
rect 4787 -1009 4833 -997
rect 4935 -121 4981 -109
rect 4935 -997 4941 -121
rect 4975 -997 4981 -121
rect 4935 -1009 4981 -997
rect 5083 -121 5129 -109
rect 5083 -997 5089 -121
rect 5123 -997 5129 -121
rect 5083 -1009 5129 -997
rect 5231 -121 5277 -109
rect 5231 -997 5237 -121
rect 5271 -997 5277 -121
rect 5231 -1009 5277 -997
rect 5379 -121 5425 -109
rect 5379 -997 5385 -121
rect 5419 -997 5425 -121
rect 5379 -1009 5425 -997
rect 5527 -121 5573 -109
rect 5527 -997 5533 -121
rect 5567 -997 5573 -121
rect 5527 -1009 5573 -997
rect -5517 -1047 -5435 -1041
rect -5517 -1081 -5505 -1047
rect -5447 -1081 -5435 -1047
rect -5517 -1087 -5435 -1081
rect -5369 -1047 -5287 -1041
rect -5369 -1081 -5357 -1047
rect -5299 -1081 -5287 -1047
rect -5369 -1087 -5287 -1081
rect -5221 -1047 -5139 -1041
rect -5221 -1081 -5209 -1047
rect -5151 -1081 -5139 -1047
rect -5221 -1087 -5139 -1081
rect -5073 -1047 -4991 -1041
rect -5073 -1081 -5061 -1047
rect -5003 -1081 -4991 -1047
rect -5073 -1087 -4991 -1081
rect -4925 -1047 -4843 -1041
rect -4925 -1081 -4913 -1047
rect -4855 -1081 -4843 -1047
rect -4925 -1087 -4843 -1081
rect -4777 -1047 -4695 -1041
rect -4777 -1081 -4765 -1047
rect -4707 -1081 -4695 -1047
rect -4777 -1087 -4695 -1081
rect -4629 -1047 -4547 -1041
rect -4629 -1081 -4617 -1047
rect -4559 -1081 -4547 -1047
rect -4629 -1087 -4547 -1081
rect -4481 -1047 -4399 -1041
rect -4481 -1081 -4469 -1047
rect -4411 -1081 -4399 -1047
rect -4481 -1087 -4399 -1081
rect -4333 -1047 -4251 -1041
rect -4333 -1081 -4321 -1047
rect -4263 -1081 -4251 -1047
rect -4333 -1087 -4251 -1081
rect -4185 -1047 -4103 -1041
rect -4185 -1081 -4173 -1047
rect -4115 -1081 -4103 -1047
rect -4185 -1087 -4103 -1081
rect -4037 -1047 -3955 -1041
rect -4037 -1081 -4025 -1047
rect -3967 -1081 -3955 -1047
rect -4037 -1087 -3955 -1081
rect -3889 -1047 -3807 -1041
rect -3889 -1081 -3877 -1047
rect -3819 -1081 -3807 -1047
rect -3889 -1087 -3807 -1081
rect -3741 -1047 -3659 -1041
rect -3741 -1081 -3729 -1047
rect -3671 -1081 -3659 -1047
rect -3741 -1087 -3659 -1081
rect -3593 -1047 -3511 -1041
rect -3593 -1081 -3581 -1047
rect -3523 -1081 -3511 -1047
rect -3593 -1087 -3511 -1081
rect -3445 -1047 -3363 -1041
rect -3445 -1081 -3433 -1047
rect -3375 -1081 -3363 -1047
rect -3445 -1087 -3363 -1081
rect -3297 -1047 -3215 -1041
rect -3297 -1081 -3285 -1047
rect -3227 -1081 -3215 -1047
rect -3297 -1087 -3215 -1081
rect -3149 -1047 -3067 -1041
rect -3149 -1081 -3137 -1047
rect -3079 -1081 -3067 -1047
rect -3149 -1087 -3067 -1081
rect -3001 -1047 -2919 -1041
rect -3001 -1081 -2989 -1047
rect -2931 -1081 -2919 -1047
rect -3001 -1087 -2919 -1081
rect -2853 -1047 -2771 -1041
rect -2853 -1081 -2841 -1047
rect -2783 -1081 -2771 -1047
rect -2853 -1087 -2771 -1081
rect -2705 -1047 -2623 -1041
rect -2705 -1081 -2693 -1047
rect -2635 -1081 -2623 -1047
rect -2705 -1087 -2623 -1081
rect -2557 -1047 -2475 -1041
rect -2557 -1081 -2545 -1047
rect -2487 -1081 -2475 -1047
rect -2557 -1087 -2475 -1081
rect -2409 -1047 -2327 -1041
rect -2409 -1081 -2397 -1047
rect -2339 -1081 -2327 -1047
rect -2409 -1087 -2327 -1081
rect -2261 -1047 -2179 -1041
rect -2261 -1081 -2249 -1047
rect -2191 -1081 -2179 -1047
rect -2261 -1087 -2179 -1081
rect -2113 -1047 -2031 -1041
rect -2113 -1081 -2101 -1047
rect -2043 -1081 -2031 -1047
rect -2113 -1087 -2031 -1081
rect -1965 -1047 -1883 -1041
rect -1965 -1081 -1953 -1047
rect -1895 -1081 -1883 -1047
rect -1965 -1087 -1883 -1081
rect -1817 -1047 -1735 -1041
rect -1817 -1081 -1805 -1047
rect -1747 -1081 -1735 -1047
rect -1817 -1087 -1735 -1081
rect -1669 -1047 -1587 -1041
rect -1669 -1081 -1657 -1047
rect -1599 -1081 -1587 -1047
rect -1669 -1087 -1587 -1081
rect -1521 -1047 -1439 -1041
rect -1521 -1081 -1509 -1047
rect -1451 -1081 -1439 -1047
rect -1521 -1087 -1439 -1081
rect -1373 -1047 -1291 -1041
rect -1373 -1081 -1361 -1047
rect -1303 -1081 -1291 -1047
rect -1373 -1087 -1291 -1081
rect -1225 -1047 -1143 -1041
rect -1225 -1081 -1213 -1047
rect -1155 -1081 -1143 -1047
rect -1225 -1087 -1143 -1081
rect -1077 -1047 -995 -1041
rect -1077 -1081 -1065 -1047
rect -1007 -1081 -995 -1047
rect -1077 -1087 -995 -1081
rect -929 -1047 -847 -1041
rect -929 -1081 -917 -1047
rect -859 -1081 -847 -1047
rect -929 -1087 -847 -1081
rect -781 -1047 -699 -1041
rect -781 -1081 -769 -1047
rect -711 -1081 -699 -1047
rect -781 -1087 -699 -1081
rect -633 -1047 -551 -1041
rect -633 -1081 -621 -1047
rect -563 -1081 -551 -1047
rect -633 -1087 -551 -1081
rect -485 -1047 -403 -1041
rect -485 -1081 -473 -1047
rect -415 -1081 -403 -1047
rect -485 -1087 -403 -1081
rect -337 -1047 -255 -1041
rect -337 -1081 -325 -1047
rect -267 -1081 -255 -1047
rect -337 -1087 -255 -1081
rect -189 -1047 -107 -1041
rect -189 -1081 -177 -1047
rect -119 -1081 -107 -1047
rect -189 -1087 -107 -1081
rect -41 -1047 41 -1041
rect -41 -1081 -29 -1047
rect 29 -1081 41 -1047
rect -41 -1087 41 -1081
rect 107 -1047 189 -1041
rect 107 -1081 119 -1047
rect 177 -1081 189 -1047
rect 107 -1087 189 -1081
rect 255 -1047 337 -1041
rect 255 -1081 267 -1047
rect 325 -1081 337 -1047
rect 255 -1087 337 -1081
rect 403 -1047 485 -1041
rect 403 -1081 415 -1047
rect 473 -1081 485 -1047
rect 403 -1087 485 -1081
rect 551 -1047 633 -1041
rect 551 -1081 563 -1047
rect 621 -1081 633 -1047
rect 551 -1087 633 -1081
rect 699 -1047 781 -1041
rect 699 -1081 711 -1047
rect 769 -1081 781 -1047
rect 699 -1087 781 -1081
rect 847 -1047 929 -1041
rect 847 -1081 859 -1047
rect 917 -1081 929 -1047
rect 847 -1087 929 -1081
rect 995 -1047 1077 -1041
rect 995 -1081 1007 -1047
rect 1065 -1081 1077 -1047
rect 995 -1087 1077 -1081
rect 1143 -1047 1225 -1041
rect 1143 -1081 1155 -1047
rect 1213 -1081 1225 -1047
rect 1143 -1087 1225 -1081
rect 1291 -1047 1373 -1041
rect 1291 -1081 1303 -1047
rect 1361 -1081 1373 -1047
rect 1291 -1087 1373 -1081
rect 1439 -1047 1521 -1041
rect 1439 -1081 1451 -1047
rect 1509 -1081 1521 -1047
rect 1439 -1087 1521 -1081
rect 1587 -1047 1669 -1041
rect 1587 -1081 1599 -1047
rect 1657 -1081 1669 -1047
rect 1587 -1087 1669 -1081
rect 1735 -1047 1817 -1041
rect 1735 -1081 1747 -1047
rect 1805 -1081 1817 -1047
rect 1735 -1087 1817 -1081
rect 1883 -1047 1965 -1041
rect 1883 -1081 1895 -1047
rect 1953 -1081 1965 -1047
rect 1883 -1087 1965 -1081
rect 2031 -1047 2113 -1041
rect 2031 -1081 2043 -1047
rect 2101 -1081 2113 -1047
rect 2031 -1087 2113 -1081
rect 2179 -1047 2261 -1041
rect 2179 -1081 2191 -1047
rect 2249 -1081 2261 -1047
rect 2179 -1087 2261 -1081
rect 2327 -1047 2409 -1041
rect 2327 -1081 2339 -1047
rect 2397 -1081 2409 -1047
rect 2327 -1087 2409 -1081
rect 2475 -1047 2557 -1041
rect 2475 -1081 2487 -1047
rect 2545 -1081 2557 -1047
rect 2475 -1087 2557 -1081
rect 2623 -1047 2705 -1041
rect 2623 -1081 2635 -1047
rect 2693 -1081 2705 -1047
rect 2623 -1087 2705 -1081
rect 2771 -1047 2853 -1041
rect 2771 -1081 2783 -1047
rect 2841 -1081 2853 -1047
rect 2771 -1087 2853 -1081
rect 2919 -1047 3001 -1041
rect 2919 -1081 2931 -1047
rect 2989 -1081 3001 -1047
rect 2919 -1087 3001 -1081
rect 3067 -1047 3149 -1041
rect 3067 -1081 3079 -1047
rect 3137 -1081 3149 -1047
rect 3067 -1087 3149 -1081
rect 3215 -1047 3297 -1041
rect 3215 -1081 3227 -1047
rect 3285 -1081 3297 -1047
rect 3215 -1087 3297 -1081
rect 3363 -1047 3445 -1041
rect 3363 -1081 3375 -1047
rect 3433 -1081 3445 -1047
rect 3363 -1087 3445 -1081
rect 3511 -1047 3593 -1041
rect 3511 -1081 3523 -1047
rect 3581 -1081 3593 -1047
rect 3511 -1087 3593 -1081
rect 3659 -1047 3741 -1041
rect 3659 -1081 3671 -1047
rect 3729 -1081 3741 -1047
rect 3659 -1087 3741 -1081
rect 3807 -1047 3889 -1041
rect 3807 -1081 3819 -1047
rect 3877 -1081 3889 -1047
rect 3807 -1087 3889 -1081
rect 3955 -1047 4037 -1041
rect 3955 -1081 3967 -1047
rect 4025 -1081 4037 -1047
rect 3955 -1087 4037 -1081
rect 4103 -1047 4185 -1041
rect 4103 -1081 4115 -1047
rect 4173 -1081 4185 -1047
rect 4103 -1087 4185 -1081
rect 4251 -1047 4333 -1041
rect 4251 -1081 4263 -1047
rect 4321 -1081 4333 -1047
rect 4251 -1087 4333 -1081
rect 4399 -1047 4481 -1041
rect 4399 -1081 4411 -1047
rect 4469 -1081 4481 -1047
rect 4399 -1087 4481 -1081
rect 4547 -1047 4629 -1041
rect 4547 -1081 4559 -1047
rect 4617 -1081 4629 -1047
rect 4547 -1087 4629 -1081
rect 4695 -1047 4777 -1041
rect 4695 -1081 4707 -1047
rect 4765 -1081 4777 -1047
rect 4695 -1087 4777 -1081
rect 4843 -1047 4925 -1041
rect 4843 -1081 4855 -1047
rect 4913 -1081 4925 -1047
rect 4843 -1087 4925 -1081
rect 4991 -1047 5073 -1041
rect 4991 -1081 5003 -1047
rect 5061 -1081 5073 -1047
rect 4991 -1087 5073 -1081
rect 5139 -1047 5221 -1041
rect 5139 -1081 5151 -1047
rect 5209 -1081 5221 -1047
rect 5139 -1087 5221 -1081
rect 5287 -1047 5369 -1041
rect 5287 -1081 5299 -1047
rect 5357 -1081 5369 -1047
rect 5287 -1087 5369 -1081
rect 5435 -1047 5517 -1041
rect 5435 -1081 5447 -1047
rect 5505 -1081 5517 -1047
rect 5435 -1087 5517 -1081
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -5664 -1166 5664 1166
string parameters w 4.5 l 0.45 m 2 nf 75 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
