magic
tech sky130A
timestamp 1663601768
<< nwell >>
rect -175 -30 605 125
<< pwell >>
rect -10 190 30 230
rect 405 195 445 235
rect -75 -345 520 -175
rect 115 -380 500 -345
<< nmos >>
rect 90 -305 105 -205
rect 180 -305 195 -205
rect 420 -305 435 -205
<< pmos >>
rect 0 0 15 100
rect 90 0 105 100
rect 330 0 345 100
rect 420 0 435 100
<< ndiff >>
rect 15 -220 90 -205
rect 15 -290 30 -220
rect 75 -290 90 -220
rect 15 -305 90 -290
rect 105 -220 180 -205
rect 105 -290 120 -220
rect 165 -290 180 -220
rect 105 -305 180 -290
rect 195 -220 270 -205
rect 345 -220 420 -205
rect 195 -290 210 -220
rect 255 -290 270 -220
rect 345 -290 360 -220
rect 405 -290 420 -220
rect 195 -305 270 -290
rect 345 -305 420 -290
rect 435 -220 510 -205
rect 435 -290 450 -220
rect 495 -290 510 -220
rect 435 -305 510 -290
<< pdiff >>
rect -75 85 0 100
rect -75 15 -60 85
rect -15 15 0 85
rect -75 0 0 15
rect 15 85 90 100
rect 15 15 30 85
rect 75 15 90 85
rect 15 0 90 15
rect 105 85 180 100
rect 255 85 330 100
rect 105 15 120 85
rect 165 15 180 85
rect 255 15 270 85
rect 315 15 330 85
rect 105 0 180 15
rect 255 0 330 15
rect 345 85 420 100
rect 345 15 360 85
rect 405 15 420 85
rect 345 0 420 15
rect 435 85 510 100
rect 435 15 450 85
rect 495 15 510 85
rect 435 0 510 15
<< ndiffc >>
rect 30 -290 75 -220
rect 120 -290 165 -220
rect 210 -290 255 -220
rect 360 -290 405 -220
rect 450 -290 495 -220
<< pdiffc >>
rect -60 15 -15 85
rect 30 15 75 85
rect 120 15 165 85
rect 270 15 315 85
rect 360 15 405 85
rect 450 15 495 85
<< psubdiff >>
rect -60 -220 15 -205
rect -60 -290 -45 -220
rect 0 -290 15 -220
rect -60 -305 15 -290
rect 270 -220 345 -205
rect 270 -290 285 -220
rect 330 -290 345 -220
rect 270 -305 345 -290
<< nsubdiff >>
rect -150 85 -75 100
rect -150 15 -135 85
rect -90 15 -75 85
rect -150 0 -75 15
rect 180 85 255 100
rect 180 15 195 85
rect 240 15 255 85
rect 180 0 255 15
rect 510 85 585 100
rect 510 15 525 85
rect 570 15 585 85
rect 510 0 585 15
<< psubdiffcont >>
rect -45 -290 0 -220
rect 285 -290 330 -220
<< nsubdiffcont >>
rect -135 15 -90 85
rect 195 15 240 85
rect 525 15 570 85
<< poly >>
rect -10 220 30 230
rect -10 195 0 220
rect 20 195 30 220
rect -10 185 30 195
rect 405 225 445 235
rect 405 200 415 225
rect 435 200 445 225
rect 405 190 445 200
rect 0 100 15 185
rect 330 165 390 175
rect 330 125 355 165
rect 385 125 390 165
rect 330 115 390 125
rect 90 100 105 115
rect 330 100 345 115
rect 420 100 435 190
rect 0 -15 15 0
rect 90 -25 105 0
rect 330 -25 345 0
rect 420 -15 435 0
rect 90 -35 145 -25
rect 90 -75 110 -35
rect 135 -75 145 -35
rect 90 -85 145 -75
rect 180 -95 220 -85
rect 180 -120 190 -95
rect 210 -120 220 -95
rect 180 -130 220 -120
rect 90 -140 130 -130
rect 90 -165 100 -140
rect 120 -165 130 -140
rect 90 -175 130 -165
rect 90 -205 105 -175
rect 180 -205 195 -130
rect 420 -205 435 -190
rect 90 -320 105 -305
rect 180 -320 195 -305
rect 420 -340 435 -305
rect 405 -350 445 -340
rect 405 -375 415 -350
rect 435 -375 445 -350
rect 405 -385 445 -375
<< polycont >>
rect 0 195 20 220
rect 415 200 435 225
rect 355 125 385 165
rect 110 -75 135 -35
rect 190 -120 210 -95
rect 100 -165 120 -140
rect 415 -375 435 -350
<< locali >>
rect -10 225 30 230
rect 405 225 445 235
rect -210 220 415 225
rect -210 200 -195 220
rect -120 200 0 220
rect -210 195 0 200
rect 20 200 415 220
rect 435 220 950 225
rect 435 200 860 220
rect 935 200 950 220
rect 20 195 950 200
rect -10 185 30 195
rect 405 190 445 195
rect 345 165 390 175
rect 345 125 355 165
rect 385 125 390 165
rect 345 115 390 125
rect -140 85 -85 95
rect -140 15 -135 85
rect -90 15 -85 85
rect -140 5 -85 15
rect -65 85 -10 95
rect -65 15 -60 85
rect -15 15 -10 85
rect -65 5 -10 15
rect 25 85 80 95
rect 25 15 30 85
rect 75 15 80 85
rect 25 0 80 15
rect 115 85 170 95
rect 115 15 120 85
rect 165 15 170 85
rect 115 5 170 15
rect 190 85 245 95
rect 190 15 195 85
rect 240 15 245 85
rect 190 5 245 15
rect 265 85 320 95
rect 265 15 270 85
rect 315 15 320 85
rect 265 5 320 15
rect 355 85 410 95
rect 355 15 360 85
rect 405 15 410 85
rect 355 0 410 15
rect 445 85 500 95
rect 445 15 450 85
rect 495 15 500 85
rect 445 5 500 15
rect 520 85 575 95
rect 520 15 525 85
rect 570 15 575 85
rect 520 5 575 15
rect 100 -35 145 -25
rect 100 -75 110 -35
rect 135 -75 145 -35
rect 100 -85 145 -75
rect 180 -95 220 -85
rect 180 -120 190 -95
rect 210 -120 220 -95
rect 180 -130 220 -120
rect 90 -140 130 -130
rect 90 -165 100 -140
rect 120 -165 130 -140
rect 90 -175 130 -165
rect -50 -220 5 -210
rect -50 -290 -45 -220
rect 0 -290 5 -220
rect -50 -300 5 -290
rect 25 -220 80 -210
rect 25 -290 30 -220
rect 75 -290 80 -220
rect 25 -300 80 -290
rect 115 -220 170 -210
rect 115 -290 120 -220
rect 165 -290 170 -220
rect 115 -300 170 -290
rect 205 -220 260 -210
rect 205 -290 210 -220
rect 255 -290 260 -220
rect 205 -300 260 -290
rect 280 -220 335 -210
rect 280 -290 285 -220
rect 330 -290 335 -220
rect 280 -300 335 -290
rect 355 -220 410 -210
rect 355 -290 360 -220
rect 405 -290 410 -220
rect 355 -300 410 -290
rect 445 -220 500 -210
rect 445 -290 450 -220
rect 495 -290 500 -220
rect 445 -300 500 -290
rect 660 -305 785 -220
rect 405 -350 445 -340
rect -210 -355 415 -350
rect -210 -375 -195 -355
rect -120 -375 415 -355
rect 435 -355 950 -350
rect 435 -375 875 -355
rect 935 -375 950 -355
rect -210 -380 950 -375
rect 405 -385 445 -380
<< viali >>
rect -200 295 940 325
rect -195 200 -120 220
rect 860 200 935 220
rect 355 125 385 165
rect -135 15 -90 85
rect -60 15 -15 85
rect 30 15 75 85
rect 120 15 165 85
rect 195 15 240 85
rect 270 15 315 85
rect 360 15 405 85
rect 450 15 495 85
rect 525 15 570 85
rect 810 15 890 55
rect 110 -75 135 -35
rect 370 -90 450 -50
rect 190 -120 210 -95
rect 100 -165 120 -140
rect -45 -290 0 -220
rect 30 -290 75 -220
rect 120 -290 165 -220
rect 210 -290 255 -220
rect 285 -290 330 -220
rect 360 -290 405 -220
rect 450 -290 495 -220
rect -195 -375 -120 -355
rect 875 -375 935 -355
rect -200 -465 935 -435
<< metal1 >>
rect -210 325 950 335
rect -210 295 -200 325
rect 940 295 950 325
rect -210 285 950 295
rect -65 230 -10 285
rect -210 220 -115 230
rect -210 200 -195 220
rect -120 200 -115 220
rect -210 190 -115 200
rect -65 185 -5 230
rect -140 85 -85 95
rect -140 15 -135 85
rect -90 15 -85 85
rect -140 5 -85 15
rect -65 85 -10 185
rect -65 15 -60 85
rect -15 15 -10 85
rect -65 5 -10 15
rect 25 85 80 95
rect 25 15 30 85
rect 75 15 80 85
rect 25 0 80 15
rect 115 85 170 285
rect 115 15 120 85
rect 165 15 170 85
rect 115 5 170 15
rect 190 85 245 285
rect 190 15 195 85
rect 240 15 245 85
rect 190 5 245 15
rect 265 85 320 285
rect 345 165 390 175
rect 345 125 355 165
rect 385 125 390 165
rect 345 115 390 125
rect 265 15 270 85
rect 315 15 320 85
rect 265 5 320 15
rect 355 85 410 95
rect 355 15 360 85
rect 405 15 410 85
rect 355 0 410 15
rect 445 85 500 285
rect 445 15 450 85
rect 495 15 500 85
rect 445 5 500 15
rect 520 85 575 285
rect 855 220 950 230
rect 855 200 860 220
rect 935 200 950 220
rect 855 190 950 200
rect 520 15 525 85
rect 570 15 575 85
rect 520 5 575 15
rect 800 55 900 65
rect 800 15 810 55
rect 890 15 900 55
rect 100 -35 145 -25
rect -210 -80 -25 -40
rect -40 -100 -25 -80
rect 100 -75 105 -35
rect 135 -75 145 -35
rect 800 -40 900 15
rect 100 -85 145 -75
rect 360 -50 950 -40
rect 180 -95 220 -85
rect 180 -100 190 -95
rect -40 -115 190 -100
rect 180 -120 190 -115
rect 210 -120 220 -95
rect 360 -90 370 -50
rect 450 -80 950 -50
rect 450 -90 460 -80
rect 360 -100 460 -90
rect 180 -130 220 -120
rect -210 -145 -25 -130
rect 90 -140 130 -130
rect 90 -145 100 -140
rect -210 -160 100 -145
rect -210 -170 -25 -160
rect 90 -165 100 -160
rect 120 -165 130 -140
rect 90 -175 130 -165
rect 610 -135 950 -130
rect 610 -165 620 -135
rect 750 -165 950 -135
rect 610 -170 950 -165
rect -50 -220 5 -210
rect -50 -290 -45 -220
rect 0 -290 5 -220
rect -210 -355 -115 -345
rect -210 -375 -195 -355
rect -120 -375 -115 -355
rect -210 -385 -115 -375
rect -50 -425 5 -290
rect 25 -220 80 -210
rect 25 -290 30 -220
rect 75 -290 80 -220
rect 25 -300 80 -290
rect 115 -220 170 -210
rect 115 -290 120 -220
rect 165 -290 170 -220
rect 115 -300 170 -290
rect 205 -220 260 -210
rect 205 -290 210 -220
rect 255 -290 260 -220
rect 205 -300 260 -290
rect 280 -220 335 -210
rect 280 -290 285 -220
rect 330 -290 335 -220
rect 280 -425 335 -290
rect 355 -220 410 -210
rect 355 -290 360 -220
rect 405 -290 410 -220
rect 355 -425 410 -290
rect 445 -220 500 -210
rect 445 -290 450 -220
rect 495 -290 500 -220
rect 445 -300 500 -290
rect 870 -355 950 -345
rect 870 -375 875 -355
rect 935 -375 950 -355
rect 870 -385 950 -375
rect -210 -435 950 -425
rect -210 -465 -200 -435
rect 935 -465 950 -435
rect -210 -475 950 -465
<< via1 >>
rect -200 295 940 325
rect -135 15 -90 85
rect 30 15 75 85
rect 355 125 385 165
rect 360 15 405 85
rect 810 15 890 55
rect 105 -75 110 -35
rect 110 -75 135 -35
rect 370 -90 450 -50
rect 620 -165 750 -135
rect 30 -290 75 -220
rect 120 -290 165 -220
rect 210 -290 255 -220
rect 450 -290 495 -220
rect -200 -465 935 -435
<< metal2 >>
rect -210 325 950 335
rect -210 295 -200 325
rect 940 295 950 325
rect -210 285 950 295
rect -140 85 -85 285
rect -140 15 -135 85
rect -90 15 -85 85
rect -140 5 -85 15
rect 25 165 665 175
rect 25 125 355 165
rect 385 125 665 165
rect 25 115 665 125
rect 25 85 80 115
rect 610 105 665 115
rect 610 95 670 105
rect 25 15 30 85
rect 75 15 80 85
rect 25 -220 80 15
rect 355 85 410 95
rect 355 15 360 85
rect 405 15 410 85
rect 355 -25 410 15
rect 95 -35 410 -25
rect 95 -75 105 -35
rect 135 -40 410 -35
rect 610 15 620 95
rect 660 15 670 95
rect 610 5 670 15
rect 800 55 900 65
rect 800 15 810 55
rect 890 15 900 55
rect 800 5 900 15
rect 135 -50 460 -40
rect 135 -75 370 -50
rect 95 -85 370 -75
rect 25 -290 30 -220
rect 75 -290 80 -220
rect 25 -300 80 -290
rect 115 -220 170 -210
rect 115 -290 120 -220
rect 165 -290 170 -220
rect 115 -325 170 -290
rect 205 -220 260 -85
rect 360 -90 370 -85
rect 450 -90 460 -50
rect 360 -100 460 -90
rect 610 -130 665 5
rect 610 -135 755 -130
rect 610 -165 620 -135
rect 750 -165 755 -135
rect 610 -170 755 -165
rect 205 -290 210 -220
rect 255 -290 260 -220
rect 205 -300 260 -290
rect 445 -220 500 -210
rect 445 -290 450 -220
rect 495 -290 500 -220
rect 445 -325 500 -290
rect 115 -380 500 -325
rect 610 -300 660 -280
rect 610 -335 620 -300
rect 650 -335 660 -300
rect 610 -425 660 -335
rect 785 -300 835 -280
rect 785 -335 795 -300
rect 825 -335 835 -300
rect 785 -425 835 -335
rect -210 -435 950 -425
rect -210 -465 -200 -435
rect 935 -465 950 -435
rect -210 -475 950 -465
<< via2 >>
rect 620 15 660 95
rect 810 15 890 55
rect 620 -335 650 -300
rect 795 -335 825 -300
rect -200 -465 935 -435
<< metal3 >>
rect 610 95 670 105
rect 610 15 620 95
rect 660 15 670 95
rect 610 5 670 15
rect 800 55 900 65
rect 800 15 810 55
rect 890 15 900 55
rect 800 5 900 15
rect 505 -300 660 -50
rect 860 -60 940 -55
rect 505 -305 620 -300
rect 610 -335 620 -305
rect 650 -335 660 -300
rect 610 -345 660 -335
rect 785 -300 940 -60
rect 785 -335 795 -300
rect 825 -305 940 -300
rect 825 -335 835 -305
rect 785 -345 835 -335
rect -210 -430 950 -425
rect -210 -465 -200 -430
rect 935 -465 950 -430
rect -210 -475 950 -465
<< via3 >>
rect 620 15 660 95
rect 810 15 890 55
rect -200 -435 935 -430
rect -200 -465 935 -435
<< mimcap >>
rect 520 -115 645 -75
rect 520 -185 550 -115
rect 620 -185 645 -115
rect 520 -275 645 -185
rect 800 -105 925 -75
rect 800 -175 815 -105
rect 885 -175 925 -105
rect 800 -275 925 -175
<< mimcapcontact >>
rect 550 -185 620 -115
rect 815 -175 885 -105
<< metal4 >>
rect 595 95 695 105
rect 595 15 620 95
rect 660 15 695 95
rect 595 -30 695 15
rect 525 -85 695 -30
rect 785 55 915 75
rect 785 15 810 55
rect 890 15 915 55
rect 530 -115 640 -85
rect 785 -95 915 15
rect 530 -185 550 -115
rect 620 -185 640 -115
rect 800 -105 900 -95
rect 800 -175 815 -105
rect 885 -175 900 -105
rect 800 -185 900 -175
rect 530 -200 640 -185
rect -210 -430 950 -425
rect -210 -465 -200 -430
rect 935 -465 950 -430
rect -210 -475 950 -465
<< labels >>
rlabel metal1 -210 -150 -210 -150 3 VIN
port 2 e
rlabel metal1 -210 -60 -210 -60 3 VIP
port 3 e
rlabel metal1 -210 210 -210 210 3 VCTRL
port 4 e
rlabel metal2 -210 310 -210 310 3 VDD
port 5 e
rlabel metal1 950 -150 950 -150 7 VOP
port 6 w
rlabel metal1 950 -60 950 -60 7 VON
port 7 w
rlabel metal1 -210 -365 -210 -365 3 PD
port 1 e
rlabel metal4 -210 -450 -210 -450 3 VSS
port 8 e
<< end >>
