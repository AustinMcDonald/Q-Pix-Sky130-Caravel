magic
tech sky130A
timestamp 1663665281
use BarePadArray  BarePadArray_0
timestamp 1663665281
transform 1 0 3195 0 1 12545
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_1
timestamp 1663665281
transform 1 0 25695 0 1 12545
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_2
timestamp 1663665281
transform 1 0 48195 0 1 12545
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_3
timestamp 1663665281
transform 1 0 70695 0 1 12545
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_4
timestamp 1663665281
transform 1 0 93195 0 1 12545
box -3080 -13385 19420 9615
<< end >>
