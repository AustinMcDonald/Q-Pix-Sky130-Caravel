magic
tech sky130A
timestamp 1663274866
use BarePadArray1x10  BarePadArray1x10_0
timestamp 1663099175
transform 1 0 -5 0 1 0
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_1
timestamp 1663099175
transform 1 0 -5 0 1 23000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_2
timestamp 1663099175
transform 1 0 -5 0 1 46000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_3
timestamp 1663099175
transform 1 0 -5 0 1 69000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_4
timestamp 1663099175
transform 1 0 -5 0 1 92000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_5
timestamp 1663099175
transform 1 0 -5 0 1 115000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_6
timestamp 1663099175
transform 1 0 -5 0 1 138000
box 0 0 225000 23000
use BarePadArray1x10  BarePadArray1x10_7
timestamp 1663099175
transform 1 0 -5 0 1 161000
box 0 0 225000 23000
<< end >>
