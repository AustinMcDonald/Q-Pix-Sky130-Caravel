magic
tech sky130A
timestamp 1663655995
<< nwell >>
rect 169142 220939 169720 220950
rect 167883 219286 169720 220939
rect 169142 219282 169720 219286
rect 189790 219288 192422 220956
rect 189790 219285 191198 219288
rect 191820 219285 192422 219288
rect 167883 196286 169720 197368
rect 169142 196282 169720 196286
rect 189790 196288 192422 197368
rect 189790 196285 191198 196288
rect 191820 196285 192422 196288
rect 167883 173286 169720 174368
rect 169142 173282 169720 173286
rect 189790 173288 192422 174368
rect 189790 173285 191198 173288
rect 191820 173285 192422 173288
rect 167883 150286 169720 151368
rect 169142 150282 169720 150286
rect 189790 150288 192422 151368
rect 189790 150285 191198 150288
rect 191820 150285 192422 150288
rect 167883 127286 169720 128368
rect 169142 127282 169720 127286
rect 189790 127288 192422 128368
rect 189790 127285 191198 127288
rect 191820 127285 192422 127288
rect 167883 104286 169720 105368
rect 169142 104282 169720 104286
rect 189790 104288 192422 105368
rect 189790 104285 191198 104288
rect 191820 104285 192422 104288
rect 167883 81286 169720 82368
rect 169142 81282 169720 81286
rect 189790 81288 192422 82368
rect 189790 81285 191198 81288
rect 191820 81285 192422 81288
rect 167883 58286 169720 59368
rect 168091 58285 168458 58286
rect 169142 58282 169720 58286
rect 189790 58288 192422 59368
rect 189790 58285 191198 58288
rect 191820 58285 192422 58288
rect 167883 35286 169720 36368
rect 169142 35282 169720 35286
rect 189790 35288 192422 36368
rect 189790 35285 191198 35288
rect 191820 35285 192422 35288
rect 167525 2357 170231 13780
rect 189044 2336 192946 13566
<< pmoslvt >>
rect 168666 220074 169466 220116
rect 190166 220074 192166 220116
rect 168666 197061 169466 197116
rect 190166 197061 192166 197116
rect 168666 174052 169466 174116
rect 190166 174052 192166 174116
rect 168666 151032 169466 151116
rect 190166 151032 192166 151116
rect 168666 128016 169466 128116
rect 190166 128016 192166 128116
rect 168666 104951 169466 105116
rect 190166 104951 192166 105116
rect 168666 81816 169466 82116
rect 190166 81816 192166 82116
rect 168666 58616 169466 59116
rect 190166 58616 192166 59116
rect 168666 35416 169466 36116
rect 190166 35416 192166 36116
rect 168666 3116 169466 13116
rect 190166 3116 192166 13116
<< pdiff >>
rect 168566 220103 168666 220116
rect 168566 220086 168578 220103
rect 168654 220086 168666 220103
rect 168566 220074 168666 220086
rect 169466 220103 169566 220116
rect 169466 220086 169478 220103
rect 169554 220086 169566 220103
rect 169466 220074 169566 220086
rect 190066 220103 190166 220116
rect 190066 220086 190078 220103
rect 190154 220086 190166 220103
rect 190066 220074 190166 220086
rect 192166 220103 192266 220116
rect 192166 220086 192178 220103
rect 192254 220086 192266 220103
rect 192166 220074 192266 220086
rect 168566 197103 168666 197116
rect 168566 197073 168578 197103
rect 168654 197073 168666 197103
rect 168566 197061 168666 197073
rect 169466 197103 169566 197116
rect 169466 197073 169478 197103
rect 169554 197073 169566 197103
rect 169466 197061 169566 197073
rect 190066 197103 190166 197116
rect 190066 197073 190078 197103
rect 190154 197073 190166 197103
rect 190066 197061 190166 197073
rect 192166 197103 192266 197116
rect 192166 197073 192178 197103
rect 192254 197073 192266 197103
rect 192166 197061 192266 197073
rect 168566 174103 168666 174116
rect 168566 174064 168578 174103
rect 168654 174064 168666 174103
rect 168566 174052 168666 174064
rect 169466 174103 169566 174116
rect 169466 174064 169478 174103
rect 169554 174064 169566 174103
rect 169466 174052 169566 174064
rect 190066 174103 190166 174116
rect 190066 174064 190078 174103
rect 190154 174064 190166 174103
rect 190066 174052 190166 174064
rect 192166 174103 192266 174116
rect 192166 174064 192178 174103
rect 192254 174064 192266 174103
rect 192166 174052 192266 174064
rect 168566 151103 168666 151116
rect 168566 151044 168578 151103
rect 168654 151044 168666 151103
rect 168566 151032 168666 151044
rect 169466 151103 169566 151116
rect 169466 151044 169478 151103
rect 169554 151044 169566 151103
rect 169466 151032 169566 151044
rect 190066 151103 190166 151116
rect 190066 151044 190078 151103
rect 190154 151044 190166 151103
rect 190066 151032 190166 151044
rect 192166 151103 192266 151116
rect 192166 151044 192178 151103
rect 192254 151044 192266 151103
rect 192166 151032 192266 151044
rect 168566 128103 168666 128116
rect 168566 128028 168578 128103
rect 168654 128028 168666 128103
rect 168566 128016 168666 128028
rect 169466 128103 169566 128116
rect 169466 128028 169478 128103
rect 169554 128028 169566 128103
rect 169466 128016 169566 128028
rect 190066 128103 190166 128116
rect 190066 128028 190078 128103
rect 190154 128028 190166 128103
rect 190066 128016 190166 128028
rect 192166 128103 192266 128116
rect 192166 128028 192178 128103
rect 192254 128028 192266 128103
rect 192166 128016 192266 128028
rect 168566 105103 168666 105116
rect 168566 104963 168578 105103
rect 168654 104963 168666 105103
rect 168566 104951 168666 104963
rect 169466 105103 169566 105116
rect 169466 104963 169478 105103
rect 169554 104963 169566 105103
rect 169466 104951 169566 104963
rect 190066 105103 190166 105116
rect 190066 104963 190078 105103
rect 190154 104963 190166 105103
rect 190066 104951 190166 104963
rect 192166 105103 192266 105116
rect 192166 104963 192178 105103
rect 192254 104963 192266 105103
rect 192166 104951 192266 104963
rect 168566 82103 168666 82116
rect 168566 81828 168578 82103
rect 168654 81828 168666 82103
rect 168566 81816 168666 81828
rect 169466 82103 169566 82116
rect 169466 81828 169478 82103
rect 169554 81828 169566 82103
rect 169466 81816 169566 81828
rect 190066 82103 190166 82116
rect 190066 81828 190078 82103
rect 190154 81828 190166 82103
rect 190066 81816 190166 81828
rect 192166 82103 192266 82116
rect 192166 81828 192178 82103
rect 192254 81828 192266 82103
rect 192166 81816 192266 81828
rect 168566 59103 168666 59116
rect 168566 58628 168578 59103
rect 168654 58628 168666 59103
rect 168566 58616 168666 58628
rect 169466 59103 169566 59116
rect 169466 58628 169478 59103
rect 169554 58628 169566 59103
rect 169466 58616 169566 58628
rect 190066 59103 190166 59116
rect 190066 58628 190078 59103
rect 190154 58628 190166 59103
rect 190066 58616 190166 58628
rect 192166 59103 192266 59116
rect 192166 58628 192178 59103
rect 192254 58628 192266 59103
rect 192166 58616 192266 58628
rect 168566 36103 168666 36116
rect 168566 35428 168578 36103
rect 168654 35428 168666 36103
rect 168566 35416 168666 35428
rect 169466 36103 169566 36116
rect 169466 35428 169478 36103
rect 169554 35428 169566 36103
rect 169466 35416 169566 35428
rect 190066 36103 190166 36116
rect 190066 35428 190078 36103
rect 190154 35428 190166 36103
rect 190066 35416 190166 35428
rect 192166 36103 192266 36116
rect 192166 35428 192178 36103
rect 192254 35428 192266 36103
rect 192166 35416 192266 35428
rect 168566 13103 168666 13116
rect 168566 3128 168578 13103
rect 168654 3128 168666 13103
rect 168566 3116 168666 3128
rect 169466 13103 169566 13116
rect 169466 3128 169478 13103
rect 169554 3128 169566 13103
rect 169466 3116 169566 3128
rect 190066 13103 190166 13116
rect 190066 3128 190078 13103
rect 190154 3128 190166 13103
rect 190066 3116 190166 3128
rect 192166 13103 192266 13116
rect 192166 3128 192178 13103
rect 192254 3128 192266 13103
rect 192166 3116 192266 3128
<< pdiffc >>
rect 168578 220086 168654 220103
rect 169478 220086 169554 220103
rect 190078 220086 190154 220103
rect 192178 220086 192254 220103
rect 168578 197073 168654 197103
rect 169478 197073 169554 197103
rect 190078 197073 190154 197103
rect 192178 197073 192254 197103
rect 168578 174064 168654 174103
rect 169478 174064 169554 174103
rect 190078 174064 190154 174103
rect 192178 174064 192254 174103
rect 168578 151044 168654 151103
rect 169478 151044 169554 151103
rect 190078 151044 190154 151103
rect 192178 151044 192254 151103
rect 168578 128028 168654 128103
rect 169478 128028 169554 128103
rect 190078 128028 190154 128103
rect 192178 128028 192254 128103
rect 168578 104963 168654 105103
rect 169478 104963 169554 105103
rect 190078 104963 190154 105103
rect 192178 104963 192254 105103
rect 168578 81828 168654 82103
rect 169478 81828 169554 82103
rect 190078 81828 190154 82103
rect 192178 81828 192254 82103
rect 168578 58628 168654 59103
rect 169478 58628 169554 59103
rect 190078 58628 190154 59103
rect 192178 58628 192254 59103
rect 168578 35428 168654 36103
rect 169478 35428 169554 36103
rect 190078 35428 190154 36103
rect 192178 35428 192254 36103
rect 168578 3128 168654 13103
rect 169478 3128 169554 13103
rect 190078 3128 190154 13103
rect 192178 3128 192254 13103
<< nsubdiff >>
rect 168466 220103 168566 220116
rect 168466 220086 168479 220103
rect 168555 220086 168566 220103
rect 168466 220074 168566 220086
rect 189966 220103 190066 220116
rect 189966 220086 189979 220103
rect 190055 220086 190066 220103
rect 189966 220074 190066 220086
rect 192266 220103 192366 220116
rect 192266 220086 192279 220103
rect 192355 220086 192366 220103
rect 192266 220074 192366 220086
rect 168466 197103 168566 197116
rect 168466 197073 168479 197103
rect 168555 197073 168566 197103
rect 168466 197061 168566 197073
rect 189966 197103 190066 197116
rect 189966 197073 189979 197103
rect 190055 197073 190066 197103
rect 189966 197061 190066 197073
rect 192266 197103 192366 197116
rect 192266 197073 192279 197103
rect 192355 197073 192366 197103
rect 192266 197061 192366 197073
rect 168466 174103 168566 174116
rect 168466 174064 168479 174103
rect 168555 174064 168566 174103
rect 168466 174052 168566 174064
rect 189966 174103 190066 174116
rect 189966 174064 189979 174103
rect 190055 174064 190066 174103
rect 189966 174052 190066 174064
rect 192266 174103 192366 174116
rect 192266 174064 192279 174103
rect 192355 174064 192366 174103
rect 192266 174052 192366 174064
rect 168466 151103 168566 151116
rect 168466 151044 168479 151103
rect 168555 151044 168566 151103
rect 168466 151032 168566 151044
rect 189966 151103 190066 151116
rect 189966 151044 189979 151103
rect 190055 151044 190066 151103
rect 189966 151032 190066 151044
rect 192266 151103 192366 151116
rect 192266 151044 192279 151103
rect 192355 151044 192366 151103
rect 192266 151032 192366 151044
rect 168466 128103 168566 128116
rect 168466 128028 168479 128103
rect 168555 128028 168566 128103
rect 168466 128016 168566 128028
rect 189966 128103 190066 128116
rect 189966 128028 189979 128103
rect 190055 128028 190066 128103
rect 189966 128016 190066 128028
rect 192266 128103 192366 128116
rect 192266 128028 192279 128103
rect 192355 128028 192366 128103
rect 192266 128016 192366 128028
rect 168466 105103 168566 105116
rect 168466 104963 168479 105103
rect 168555 104963 168566 105103
rect 168466 104951 168566 104963
rect 189966 105103 190066 105116
rect 189966 104963 189979 105103
rect 190055 104963 190066 105103
rect 189966 104951 190066 104963
rect 192266 105103 192366 105116
rect 192266 104963 192279 105103
rect 192355 104963 192366 105103
rect 192266 104951 192366 104963
rect 168466 82103 168566 82116
rect 168466 81828 168479 82103
rect 168555 81828 168566 82103
rect 168466 81816 168566 81828
rect 189966 82103 190066 82116
rect 189966 81828 189979 82103
rect 190055 81828 190066 82103
rect 189966 81816 190066 81828
rect 192266 82103 192366 82116
rect 192266 81828 192279 82103
rect 192355 81828 192366 82103
rect 192266 81816 192366 81828
rect 168466 59103 168566 59116
rect 168466 58628 168479 59103
rect 168555 58628 168566 59103
rect 168466 58616 168566 58628
rect 189966 59103 190066 59116
rect 189966 58628 189979 59103
rect 190055 58628 190066 59103
rect 189966 58616 190066 58628
rect 192266 59103 192366 59116
rect 192266 58628 192279 59103
rect 192355 58628 192366 59103
rect 192266 58616 192366 58628
rect 168466 36103 168566 36116
rect 168466 35428 168479 36103
rect 168555 35428 168566 36103
rect 168466 35416 168566 35428
rect 189966 36103 190066 36116
rect 189966 35428 189979 36103
rect 190055 35428 190066 36103
rect 189966 35416 190066 35428
rect 192266 36103 192366 36116
rect 192266 35428 192279 36103
rect 192355 35428 192366 36103
rect 192266 35416 192366 35428
rect 168466 13103 168566 13116
rect 168466 3128 168479 13103
rect 168555 3128 168566 13103
rect 168466 3116 168566 3128
rect 189966 13103 190066 13116
rect 189966 3128 189979 13103
rect 190055 3128 190066 13103
rect 189966 3116 190066 3128
rect 192266 13103 192366 13116
rect 192266 3128 192279 13103
rect 192355 3128 192366 13103
rect 192266 3116 192366 3128
<< nsubdiffcont >>
rect 168479 220086 168555 220103
rect 189979 220086 190055 220103
rect 192279 220086 192355 220103
rect 168479 197073 168555 197103
rect 189979 197073 190055 197103
rect 192279 197073 192355 197103
rect 168479 174064 168555 174103
rect 189979 174064 190055 174103
rect 192279 174064 192355 174103
rect 168479 151044 168555 151103
rect 189979 151044 190055 151103
rect 192279 151044 192355 151103
rect 168479 128028 168555 128103
rect 189979 128028 190055 128103
rect 192279 128028 192355 128103
rect 168479 104963 168555 105103
rect 189979 104963 190055 105103
rect 192279 104963 192355 105103
rect 168479 81828 168555 82103
rect 189979 81828 190055 82103
rect 192279 81828 192355 82103
rect 168479 58628 168555 59103
rect 189979 58628 190055 59103
rect 192279 58628 192355 59103
rect 168479 35428 168555 36103
rect 189979 35428 190055 36103
rect 192279 35428 192355 36103
rect 168479 3128 168555 13103
rect 189979 3128 190055 13103
rect 192279 3128 192355 13103
<< poly >>
rect 168649 220183 169462 220191
rect 168649 220149 168657 220183
rect 168649 220148 168680 220149
rect 169445 220148 169462 220183
rect 168649 220141 169462 220148
rect 190171 220184 192155 220191
rect 190171 220150 190186 220184
rect 192127 220150 192155 220184
rect 190171 220149 191157 220150
rect 191191 220149 192155 220150
rect 190171 220141 192155 220149
rect 168666 220116 169466 220141
rect 190166 220116 192166 220141
rect 168666 220059 169466 220074
rect 190166 220059 192166 220074
rect 168649 197183 169462 197191
rect 168649 197149 168657 197183
rect 168649 197148 168680 197149
rect 169445 197148 169462 197183
rect 168649 197141 169462 197148
rect 190171 197184 192155 197191
rect 190171 197150 190186 197184
rect 192127 197150 192155 197184
rect 190171 197149 191157 197150
rect 191191 197149 192155 197150
rect 190171 197141 192155 197149
rect 168666 197116 169466 197141
rect 190166 197116 192166 197141
rect 168666 197048 169466 197061
rect 190166 197048 192166 197061
rect 168649 174183 169462 174191
rect 168649 174149 168657 174183
rect 168649 174148 168680 174149
rect 169445 174148 169462 174183
rect 168649 174141 169462 174148
rect 190171 174184 192155 174191
rect 190171 174150 190186 174184
rect 192127 174150 192155 174184
rect 190171 174149 191157 174150
rect 191191 174149 192155 174150
rect 190171 174141 192155 174149
rect 168666 174116 169466 174141
rect 190166 174116 192166 174141
rect 168666 174039 169466 174052
rect 190166 174039 192166 174052
rect 168649 151183 169462 151191
rect 168649 151149 168657 151183
rect 168649 151148 168680 151149
rect 169445 151148 169462 151183
rect 168649 151141 169462 151148
rect 190171 151184 192155 151191
rect 190171 151150 190186 151184
rect 192127 151150 192155 151184
rect 190171 151149 191157 151150
rect 191191 151149 192155 151150
rect 190171 151141 192155 151149
rect 168666 151116 169466 151141
rect 190166 151116 192166 151141
rect 168666 151012 169466 151032
rect 190166 151012 192166 151032
rect 168649 128183 169462 128191
rect 168649 128149 168657 128183
rect 168649 128148 168680 128149
rect 169445 128148 169462 128183
rect 168649 128141 169462 128148
rect 190171 128184 192155 128191
rect 190171 128150 190186 128184
rect 192127 128150 192155 128184
rect 190171 128149 191157 128150
rect 191191 128149 192155 128150
rect 190171 128141 192155 128149
rect 168666 128116 169466 128141
rect 190166 128116 192166 128141
rect 168666 127987 169466 128016
rect 190166 127986 192166 128016
rect 168649 105183 169462 105191
rect 168649 105149 168657 105183
rect 168649 105148 168680 105149
rect 169445 105148 169462 105183
rect 168649 105141 169462 105148
rect 190171 105184 192155 105191
rect 190171 105150 190186 105184
rect 192127 105150 192155 105184
rect 190171 105149 191157 105150
rect 191191 105149 192155 105150
rect 190171 105141 192155 105149
rect 168666 105116 169466 105141
rect 190166 105116 192166 105141
rect 168666 104929 169466 104951
rect 190166 104935 192166 104951
rect 168649 82183 169462 82191
rect 168649 82149 168657 82183
rect 168649 82148 168680 82149
rect 169445 82148 169462 82183
rect 168649 82141 169462 82148
rect 190171 82184 192155 82191
rect 190171 82150 190186 82184
rect 192127 82150 192155 82184
rect 190171 82149 191157 82150
rect 191191 82149 192155 82150
rect 190171 82141 192155 82149
rect 168666 82116 169466 82141
rect 190166 82116 192166 82141
rect 168666 81797 169466 81816
rect 190166 81795 192166 81816
rect 168649 59183 169462 59191
rect 168649 59149 168657 59183
rect 168649 59148 168680 59149
rect 169445 59148 169462 59183
rect 168649 59141 169462 59148
rect 190171 59184 192155 59191
rect 190171 59150 190186 59184
rect 192127 59150 192155 59184
rect 190171 59149 191157 59150
rect 191191 59149 192155 59150
rect 190171 59141 192155 59149
rect 168666 59116 169466 59141
rect 190166 59116 192166 59141
rect 168666 58598 169466 58616
rect 190166 58545 192166 58616
rect 168649 36183 169462 36191
rect 168649 36149 168657 36183
rect 168649 36148 168680 36149
rect 169445 36148 169462 36183
rect 168649 36141 169462 36148
rect 190171 36184 192155 36191
rect 190171 36150 190186 36184
rect 192127 36150 192155 36184
rect 190171 36149 191157 36150
rect 191191 36149 192155 36150
rect 190171 36141 192155 36149
rect 168666 36116 169466 36141
rect 190166 36116 192166 36141
rect 168666 35388 169466 35416
rect 190166 35399 192166 35416
rect 168649 13183 169462 13191
rect 168649 13149 168657 13183
rect 168649 13148 168680 13149
rect 169445 13148 169462 13183
rect 168649 13141 169462 13148
rect 190171 13184 192155 13191
rect 190171 13150 190186 13184
rect 192127 13150 192155 13184
rect 190171 13149 191157 13150
rect 191191 13149 192155 13150
rect 190171 13141 192155 13149
rect 168666 13116 169466 13141
rect 190166 13116 192166 13141
rect 168666 3091 169466 3116
rect 190166 3092 192166 3116
<< polycont >>
rect 168657 220149 169445 220183
rect 168680 220148 169445 220149
rect 190186 220150 192127 220184
rect 191157 220149 191191 220150
rect 168657 197149 169445 197183
rect 168680 197148 169445 197149
rect 190186 197150 192127 197184
rect 191157 197149 191191 197150
rect 168657 174149 169445 174183
rect 168680 174148 169445 174149
rect 190186 174150 192127 174184
rect 191157 174149 191191 174150
rect 168657 151149 169445 151183
rect 168680 151148 169445 151149
rect 190186 151150 192127 151184
rect 191157 151149 191191 151150
rect 168657 128149 169445 128183
rect 168680 128148 169445 128149
rect 190186 128150 192127 128184
rect 191157 128149 191191 128150
rect 168657 105149 169445 105183
rect 168680 105148 169445 105149
rect 190186 105150 192127 105184
rect 191157 105149 191191 105150
rect 168657 82149 169445 82183
rect 168680 82148 169445 82149
rect 190186 82150 192127 82184
rect 191157 82149 191191 82150
rect 168657 59149 169445 59183
rect 168680 59148 169445 59149
rect 190186 59150 192127 59184
rect 191157 59149 191191 59150
rect 168657 36149 169445 36183
rect 168680 36148 169445 36149
rect 190186 36150 192127 36184
rect 191157 36149 191191 36150
rect 168657 13149 169445 13183
rect 168680 13148 169445 13149
rect 190186 13150 192127 13184
rect 191157 13149 191191 13150
<< locali >>
rect 168649 220183 169463 220191
rect 168649 220149 168657 220183
rect 168649 220148 168680 220149
rect 169445 220148 169463 220183
rect 168649 220141 169463 220148
rect 190176 220184 192154 220191
rect 190176 220150 190186 220184
rect 192127 220150 192154 220184
rect 190176 220149 191157 220150
rect 191191 220149 192154 220150
rect 190176 220146 192154 220149
rect 191149 220141 191199 220146
rect 168468 220103 168556 220114
rect 168468 220086 168474 220103
rect 168555 220086 168556 220103
rect 168468 220076 168556 220086
rect 168576 220103 168664 220114
rect 168576 220086 168578 220103
rect 168654 220086 168664 220103
rect 168576 220076 168664 220086
rect 169468 220103 169564 220114
rect 169468 220086 169478 220103
rect 169559 220086 169564 220103
rect 169468 220076 169564 220086
rect 189968 220103 190056 220114
rect 189968 220086 189974 220103
rect 190055 220086 190056 220103
rect 189968 220076 190056 220086
rect 190076 220103 190164 220114
rect 190076 220086 190078 220103
rect 190154 220086 190164 220103
rect 190076 220076 190164 220086
rect 192168 220103 192356 220114
rect 192168 220086 192178 220103
rect 192259 220086 192279 220103
rect 192355 220086 192356 220103
rect 192168 220076 192356 220086
rect 168649 197183 169463 197191
rect 168649 197149 168657 197183
rect 168649 197148 168680 197149
rect 169445 197148 169463 197183
rect 168649 197141 169463 197148
rect 190176 197184 192154 197191
rect 190176 197150 190186 197184
rect 192127 197150 192154 197184
rect 190176 197149 191157 197150
rect 191191 197149 192154 197150
rect 190176 197146 192154 197149
rect 191149 197141 191199 197146
rect 168468 197103 168556 197114
rect 168468 197073 168474 197103
rect 168555 197073 168556 197103
rect 168468 197063 168556 197073
rect 168576 197103 168664 197114
rect 168576 197073 168578 197103
rect 168654 197073 168664 197103
rect 168576 197063 168664 197073
rect 169468 197103 169564 197114
rect 169468 197073 169478 197103
rect 169559 197073 169564 197103
rect 169468 197063 169564 197073
rect 189968 197103 190056 197114
rect 189968 197073 189974 197103
rect 190055 197073 190056 197103
rect 189968 197063 190056 197073
rect 190076 197103 190164 197114
rect 190076 197073 190078 197103
rect 190154 197073 190164 197103
rect 190076 197063 190164 197073
rect 192168 197103 192356 197114
rect 192168 197073 192178 197103
rect 192259 197073 192279 197103
rect 192355 197073 192356 197103
rect 192168 197063 192356 197073
rect 168649 174183 169463 174191
rect 168649 174149 168657 174183
rect 168649 174148 168680 174149
rect 169445 174148 169463 174183
rect 168649 174141 169463 174148
rect 190176 174184 192154 174191
rect 190176 174150 190186 174184
rect 192127 174150 192154 174184
rect 190176 174149 191157 174150
rect 191191 174149 192154 174150
rect 190176 174146 192154 174149
rect 191149 174141 191199 174146
rect 168468 174103 168556 174114
rect 168468 174064 168474 174103
rect 168555 174064 168556 174103
rect 168468 174054 168556 174064
rect 168576 174103 168664 174114
rect 168576 174064 168578 174103
rect 168654 174064 168664 174103
rect 168576 174054 168664 174064
rect 169468 174103 169564 174114
rect 169468 174064 169478 174103
rect 169559 174064 169564 174103
rect 169468 174054 169564 174064
rect 189968 174103 190056 174114
rect 189968 174064 189974 174103
rect 190055 174064 190056 174103
rect 189968 174054 190056 174064
rect 190076 174103 190164 174114
rect 190076 174064 190078 174103
rect 190154 174064 190164 174103
rect 190076 174054 190164 174064
rect 192168 174103 192356 174114
rect 192168 174064 192178 174103
rect 192259 174064 192279 174103
rect 192355 174064 192356 174103
rect 192168 174054 192356 174064
rect 168649 151183 169463 151191
rect 168649 151149 168657 151183
rect 168649 151148 168680 151149
rect 169445 151148 169463 151183
rect 168649 151141 169463 151148
rect 190176 151184 192154 151191
rect 190176 151150 190186 151184
rect 192127 151150 192154 151184
rect 190176 151149 191157 151150
rect 191191 151149 192154 151150
rect 190176 151146 192154 151149
rect 191149 151141 191199 151146
rect 168468 151103 168556 151114
rect 168468 151044 168474 151103
rect 168555 151044 168556 151103
rect 168468 151034 168556 151044
rect 168576 151103 168664 151114
rect 168576 151044 168578 151103
rect 168654 151044 168664 151103
rect 168576 151034 168664 151044
rect 169468 151103 169564 151114
rect 169468 151044 169478 151103
rect 169559 151044 169564 151103
rect 169468 151034 169564 151044
rect 189968 151103 190056 151114
rect 189968 151044 189974 151103
rect 190055 151044 190056 151103
rect 189968 151034 190056 151044
rect 190076 151103 190164 151114
rect 190076 151044 190078 151103
rect 190154 151044 190164 151103
rect 190076 151034 190164 151044
rect 192168 151103 192356 151114
rect 192168 151044 192178 151103
rect 192259 151044 192279 151103
rect 192355 151044 192356 151103
rect 192168 151034 192356 151044
rect 168649 128183 169463 128191
rect 168649 128149 168657 128183
rect 168649 128148 168680 128149
rect 169445 128148 169463 128183
rect 168649 128141 169463 128148
rect 190176 128184 192154 128191
rect 190176 128150 190186 128184
rect 192127 128150 192154 128184
rect 190176 128149 191157 128150
rect 191191 128149 192154 128150
rect 190176 128146 192154 128149
rect 191149 128141 191199 128146
rect 168468 128103 168556 128114
rect 168468 128028 168474 128103
rect 168555 128028 168556 128103
rect 168468 128018 168556 128028
rect 168576 128103 168664 128114
rect 168576 128028 168578 128103
rect 168654 128028 168664 128103
rect 168576 128018 168664 128028
rect 169468 128103 169564 128114
rect 169468 128028 169478 128103
rect 169559 128028 169564 128103
rect 169468 128018 169564 128028
rect 189968 128103 190056 128114
rect 189968 128028 189974 128103
rect 190055 128028 190056 128103
rect 189968 128018 190056 128028
rect 190076 128103 190164 128114
rect 190076 128028 190078 128103
rect 190154 128028 190164 128103
rect 190076 128018 190164 128028
rect 192168 128103 192356 128114
rect 192168 128028 192178 128103
rect 192259 128028 192279 128103
rect 192355 128028 192356 128103
rect 192168 128018 192356 128028
rect 168649 105183 169463 105191
rect 168649 105149 168657 105183
rect 168649 105148 168680 105149
rect 169445 105148 169463 105183
rect 168649 105141 169463 105148
rect 190176 105184 192154 105191
rect 190176 105150 190186 105184
rect 192127 105150 192154 105184
rect 190176 105149 191157 105150
rect 191191 105149 192154 105150
rect 190176 105146 192154 105149
rect 191149 105141 191199 105146
rect 168468 105103 168556 105114
rect 168468 104963 168474 105103
rect 168555 104963 168556 105103
rect 168468 104953 168556 104963
rect 168576 105103 168664 105114
rect 168576 104963 168578 105103
rect 168654 104963 168664 105103
rect 168576 104953 168664 104963
rect 169468 105103 169564 105114
rect 169468 104963 169478 105103
rect 169559 104963 169564 105103
rect 169468 104953 169564 104963
rect 189968 105103 190056 105114
rect 189968 104963 189974 105103
rect 190055 104963 190056 105103
rect 189968 104953 190056 104963
rect 190076 105103 190164 105114
rect 190076 104963 190078 105103
rect 190154 104963 190164 105103
rect 190076 104953 190164 104963
rect 192168 105103 192356 105114
rect 192168 104963 192178 105103
rect 192259 104963 192279 105103
rect 192355 104963 192356 105103
rect 192168 104953 192356 104963
rect 168649 82183 169463 82191
rect 168649 82149 168657 82183
rect 168649 82148 168680 82149
rect 169445 82148 169463 82183
rect 168649 82141 169463 82148
rect 190176 82184 192154 82191
rect 190176 82150 190186 82184
rect 192127 82150 192154 82184
rect 190176 82149 191157 82150
rect 191191 82149 192154 82150
rect 190176 82146 192154 82149
rect 191149 82141 191199 82146
rect 168468 82103 168556 82114
rect 168468 81828 168474 82103
rect 168555 81828 168556 82103
rect 168468 81818 168556 81828
rect 168576 82103 168664 82114
rect 168576 81828 168578 82103
rect 168654 81828 168664 82103
rect 168576 81818 168664 81828
rect 169468 82103 169564 82114
rect 169468 81828 169478 82103
rect 169559 81828 169564 82103
rect 169468 81818 169564 81828
rect 189968 82103 190056 82114
rect 189968 81828 189974 82103
rect 190055 81828 190056 82103
rect 189968 81818 190056 81828
rect 190076 82103 190164 82114
rect 190076 81828 190078 82103
rect 190154 81828 190164 82103
rect 190076 81818 190164 81828
rect 192168 82103 192356 82114
rect 192168 81828 192178 82103
rect 192259 81828 192279 82103
rect 192355 81828 192356 82103
rect 192168 81818 192356 81828
rect 168649 59183 169463 59191
rect 168649 59149 168657 59183
rect 168649 59148 168680 59149
rect 169445 59148 169463 59183
rect 168649 59141 169463 59148
rect 190176 59184 192154 59191
rect 190176 59150 190186 59184
rect 192127 59150 192154 59184
rect 190176 59149 191157 59150
rect 191191 59149 192154 59150
rect 190176 59146 192154 59149
rect 191149 59141 191199 59146
rect 168468 59103 168556 59114
rect 168468 58628 168474 59103
rect 168555 58628 168556 59103
rect 168468 58618 168556 58628
rect 168576 59103 168664 59114
rect 168576 58628 168578 59103
rect 168654 58628 168664 59103
rect 168576 58618 168664 58628
rect 169468 59103 169564 59114
rect 169468 58628 169478 59103
rect 169559 58628 169564 59103
rect 169468 58618 169564 58628
rect 189968 59103 190056 59114
rect 189968 58628 189974 59103
rect 190055 58628 190056 59103
rect 189968 58618 190056 58628
rect 190076 59103 190164 59114
rect 190076 58628 190078 59103
rect 190154 58628 190164 59103
rect 190076 58618 190164 58628
rect 192168 59103 192356 59114
rect 192168 58628 192178 59103
rect 192259 58628 192279 59103
rect 192355 58628 192356 59103
rect 192168 58618 192356 58628
rect 168649 36183 169463 36191
rect 168649 36149 168657 36183
rect 168649 36148 168680 36149
rect 169445 36148 169463 36183
rect 168649 36141 169463 36148
rect 190176 36184 192154 36191
rect 190176 36150 190186 36184
rect 192127 36150 192154 36184
rect 190176 36149 191157 36150
rect 191191 36149 192154 36150
rect 190176 36146 192154 36149
rect 191149 36141 191199 36146
rect 168468 36103 168556 36114
rect 168468 35428 168474 36103
rect 168555 35428 168556 36103
rect 168468 35418 168556 35428
rect 168576 36103 168664 36114
rect 168576 35428 168578 36103
rect 168654 35428 168664 36103
rect 168576 35418 168664 35428
rect 169468 36103 169564 36114
rect 169468 35428 169478 36103
rect 169559 35428 169564 36103
rect 169468 35418 169564 35428
rect 189968 36103 190056 36114
rect 189968 35428 189974 36103
rect 190055 35428 190056 36103
rect 189968 35418 190056 35428
rect 190076 36103 190164 36114
rect 190076 35428 190078 36103
rect 190154 35428 190164 36103
rect 190076 35418 190164 35428
rect 192168 36103 192356 36114
rect 192168 35428 192178 36103
rect 192259 35428 192279 36103
rect 192355 35428 192356 36103
rect 192168 35418 192356 35428
rect 168649 13183 169463 13191
rect 168649 13149 168657 13183
rect 168649 13148 168680 13149
rect 169445 13148 169463 13183
rect 168649 13141 169463 13148
rect 190176 13184 192154 13191
rect 190176 13150 190186 13184
rect 192127 13150 192154 13184
rect 190176 13149 191157 13150
rect 191191 13149 192154 13150
rect 190176 13146 192154 13149
rect 191149 13141 191199 13146
rect 168468 13103 168556 13114
rect 168468 3128 168474 13103
rect 168555 3128 168556 13103
rect 168468 3118 168556 3128
rect 168576 13103 168664 13114
rect 168576 3128 168578 13103
rect 168654 3128 168664 13103
rect 168576 3118 168664 3128
rect 169468 13103 169564 13114
rect 169468 3128 169478 13103
rect 169559 3128 169564 13103
rect 169468 3118 169564 3128
rect 189968 13103 190056 13114
rect 189968 3128 189974 13103
rect 190055 3128 190056 13103
rect 189968 3118 190056 3128
rect 190076 13103 190164 13114
rect 190076 3128 190078 13103
rect 190154 3128 190164 13103
rect 190076 3118 190164 3128
rect 192168 13103 192356 13114
rect 192168 3128 192178 13103
rect 192259 3128 192279 13103
rect 192355 3128 192356 13103
rect 192168 3118 192356 3128
<< viali >>
rect 168657 220150 169445 220183
rect 168680 220148 169445 220150
rect 190186 220150 192127 220184
rect 168474 220086 168479 220103
rect 168479 220086 168538 220103
rect 168583 220086 168647 220103
rect 169484 220086 169554 220103
rect 169554 220086 169559 220103
rect 189974 220086 189979 220103
rect 189979 220086 190038 220103
rect 190083 220086 190147 220103
rect 192184 220086 192254 220103
rect 192254 220086 192259 220103
rect 168657 197150 169445 197183
rect 168680 197148 169445 197150
rect 190186 197150 192127 197184
rect 168474 197073 168479 197103
rect 168479 197073 168538 197103
rect 168583 197073 168647 197103
rect 169484 197073 169554 197103
rect 169554 197073 169559 197103
rect 189974 197073 189979 197103
rect 189979 197073 190038 197103
rect 190083 197073 190147 197103
rect 192184 197073 192254 197103
rect 192254 197073 192259 197103
rect 168657 174150 169445 174183
rect 168680 174148 169445 174150
rect 190186 174150 192127 174184
rect 168474 174064 168479 174103
rect 168479 174064 168538 174103
rect 168583 174064 168647 174103
rect 169484 174064 169554 174103
rect 169554 174064 169559 174103
rect 189974 174064 189979 174103
rect 189979 174064 190038 174103
rect 190083 174064 190147 174103
rect 192184 174064 192254 174103
rect 192254 174064 192259 174103
rect 168657 151150 169445 151183
rect 168680 151148 169445 151150
rect 190186 151150 192127 151184
rect 168474 151044 168479 151103
rect 168479 151044 168538 151103
rect 168583 151044 168647 151103
rect 169484 151044 169554 151103
rect 169554 151044 169559 151103
rect 189974 151044 189979 151103
rect 189979 151044 190038 151103
rect 190083 151044 190147 151103
rect 192184 151044 192254 151103
rect 192254 151044 192259 151103
rect 168657 128150 169445 128183
rect 168680 128148 169445 128150
rect 190186 128150 192127 128184
rect 168474 128028 168479 128103
rect 168479 128028 168538 128103
rect 168583 128028 168647 128103
rect 169484 128028 169554 128103
rect 169554 128028 169559 128103
rect 189974 128028 189979 128103
rect 189979 128028 190038 128103
rect 190083 128028 190147 128103
rect 192184 128028 192254 128103
rect 192254 128028 192259 128103
rect 168657 105150 169445 105183
rect 168680 105148 169445 105150
rect 190186 105150 192127 105184
rect 168474 104963 168479 105103
rect 168479 104963 168538 105103
rect 168583 104963 168647 105103
rect 169484 104963 169554 105103
rect 169554 104963 169559 105103
rect 189974 104963 189979 105103
rect 189979 104963 190038 105103
rect 190083 104963 190147 105103
rect 192184 104963 192254 105103
rect 192254 104963 192259 105103
rect 168657 82150 169445 82183
rect 168680 82148 169445 82150
rect 190186 82150 192127 82184
rect 168474 81828 168479 82103
rect 168479 81828 168538 82103
rect 168583 81828 168647 82103
rect 169484 81828 169554 82103
rect 169554 81828 169559 82103
rect 189974 81828 189979 82103
rect 189979 81828 190038 82103
rect 190083 81828 190147 82103
rect 192184 81828 192254 82103
rect 192254 81828 192259 82103
rect 168657 59150 169445 59183
rect 168680 59148 169445 59150
rect 190186 59150 192127 59184
rect 168474 58628 168479 59103
rect 168479 58628 168538 59103
rect 168583 58628 168647 59103
rect 169484 58628 169554 59103
rect 169554 58628 169559 59103
rect 189974 58628 189979 59103
rect 189979 58628 190038 59103
rect 190083 58628 190147 59103
rect 192184 58628 192254 59103
rect 192254 58628 192259 59103
rect 168657 36150 169445 36183
rect 168680 36148 169445 36150
rect 190186 36150 192127 36184
rect 168474 35428 168479 36103
rect 168479 35428 168538 36103
rect 168583 35428 168647 36103
rect 169484 35428 169554 36103
rect 169554 35428 169559 36103
rect 189974 35428 189979 36103
rect 189979 35428 190038 36103
rect 190083 35428 190147 36103
rect 192184 35428 192254 36103
rect 192254 35428 192259 36103
rect 168657 13150 169445 13183
rect 168680 13148 169445 13150
rect 190186 13150 192127 13184
rect 168474 3128 168479 13103
rect 168479 3128 168538 13103
rect 168583 3128 168647 13103
rect 169484 3128 169554 13103
rect 169554 3128 169559 13103
rect 189974 3128 189979 13103
rect 189979 3128 190038 13103
rect 190083 3128 190147 13103
rect 192184 3128 192254 13103
rect 192254 3128 192259 13103
<< metal1 >>
rect 167245 220515 168745 221020
rect 189745 220736 191245 221020
rect 189745 220515 190941 220736
rect 191091 220515 191245 220736
rect 168468 220307 168545 220515
rect 168468 220103 168546 220307
rect 168649 220183 170535 220203
rect 168649 220150 168657 220183
rect 168649 220148 168680 220150
rect 169445 220148 170535 220183
rect 168649 220141 170535 220148
rect 189967 220120 190046 220515
rect 192749 220203 193020 220204
rect 190171 220184 193020 220203
rect 190171 220150 190186 220184
rect 192127 220150 193020 220184
rect 190171 220141 193020 220150
rect 190171 220137 192166 220141
rect 168468 220086 168474 220103
rect 168538 220086 168546 220103
rect 168468 220077 168546 220086
rect 168576 220103 168654 220113
rect 168576 220086 168583 220103
rect 168647 220086 168654 220103
rect 168576 219916 168654 220086
rect 169478 220103 169566 220114
rect 169478 220086 169484 220103
rect 169559 220086 169566 220103
rect 169478 220059 169566 220086
rect 189968 220103 190046 220120
rect 189968 220086 189974 220103
rect 190038 220086 190046 220103
rect 189968 220077 190046 220086
rect 190076 220103 190154 220113
rect 190076 220086 190083 220103
rect 190147 220086 190154 220103
rect 168575 219896 168654 219916
rect 169480 219896 169566 220059
rect 190076 219916 190154 220086
rect 192178 220103 192266 220114
rect 192178 220086 192184 220103
rect 192259 220086 192266 220103
rect 192178 220066 192266 220086
rect 190075 219896 190154 219916
rect 168575 219839 168653 219896
rect 168373 219771 168653 219839
rect 166480 219762 166985 219764
rect 168373 219763 168652 219771
rect 167708 219762 168652 219763
rect 166480 219728 168652 219762
rect 166480 219321 168449 219728
rect 168574 219725 168652 219728
rect 166480 219320 167724 219321
rect 166480 218244 166985 219320
rect 167245 219319 167724 219320
rect 169435 216392 169912 219896
rect 190075 219869 190153 219896
rect 189429 219867 190153 219869
rect 188985 219734 190153 219867
rect 192177 219824 192266 220066
rect 192177 219797 192267 219824
rect 188985 218027 189484 219734
rect 190075 219733 190153 219734
rect 192178 219606 192267 219797
rect 192177 219555 192267 219606
rect 192177 219132 192266 219555
rect 192177 219107 192267 219132
rect 192178 218904 192267 219107
rect 192104 216333 192426 218904
rect 168223 197357 168724 197817
rect 168468 197307 168545 197357
rect 168468 197103 168546 197307
rect 170510 197203 171015 197368
rect 189837 197367 190147 197928
rect 168649 197183 171015 197203
rect 168649 197150 168657 197183
rect 168649 197148 168680 197150
rect 169445 197148 171015 197183
rect 168649 197141 171015 197148
rect 168468 197073 168474 197103
rect 168538 197073 168546 197103
rect 168468 197064 168546 197073
rect 168576 197103 168654 197113
rect 168576 197073 168583 197103
rect 168647 197073 168654 197103
rect 168576 196916 168654 197073
rect 169478 197103 169566 197114
rect 169478 197073 169484 197103
rect 169559 197073 169566 197103
rect 169478 197059 169566 197073
rect 168575 196896 168654 196916
rect 169480 196896 169566 197059
rect 168575 196839 168653 196896
rect 168373 196771 168653 196839
rect 166480 196762 166985 196764
rect 168373 196763 168652 196771
rect 167708 196762 168652 196763
rect 166480 196728 168652 196762
rect 166480 196321 168449 196728
rect 168574 196725 168652 196728
rect 166480 196320 167724 196321
rect 166480 193650 166985 196320
rect 167245 196319 167724 196320
rect 169435 193791 169912 196896
rect 170510 195755 171015 197141
rect 189967 197120 190046 197367
rect 193010 197204 193515 197368
rect 192749 197203 193515 197204
rect 190171 197184 193515 197203
rect 190171 197150 190186 197184
rect 192127 197150 193515 197184
rect 190171 197141 193515 197150
rect 190171 197137 192166 197141
rect 189968 197103 190046 197120
rect 189968 197073 189974 197103
rect 190038 197073 190046 197103
rect 189968 197064 190046 197073
rect 190076 197103 190154 197113
rect 190076 197073 190083 197103
rect 190147 197073 190154 197103
rect 190076 196916 190154 197073
rect 192178 197103 192266 197114
rect 192178 197073 192184 197103
rect 192259 197073 192266 197103
rect 192178 197066 192266 197073
rect 190075 196896 190154 196916
rect 190075 196869 190153 196896
rect 189429 196867 190153 196869
rect 188985 196734 190153 196867
rect 192177 196824 192266 197066
rect 192177 196797 192267 196824
rect 188985 195250 189484 196734
rect 190075 196733 190153 196734
rect 192178 196606 192267 196797
rect 192177 196555 192267 196606
rect 192177 196132 192266 196555
rect 192177 196107 192267 196132
rect 192178 195904 192267 196107
rect 169418 193331 169919 193791
rect 188980 193650 189485 195250
rect 192104 194023 192426 195904
rect 193010 195755 193515 197141
rect 192104 193650 192427 194023
rect 192109 193266 192427 193650
rect 168286 174827 168734 174832
rect 168280 174372 168734 174827
rect 168280 174367 168728 174372
rect 189764 174368 190212 174828
rect 168468 174307 168545 174367
rect 168468 174103 168546 174307
rect 170510 174203 171015 174368
rect 168649 174183 171015 174203
rect 168649 174150 168657 174183
rect 168649 174148 168680 174150
rect 169445 174148 171015 174183
rect 168649 174141 171015 174148
rect 168468 174064 168474 174103
rect 168538 174064 168546 174103
rect 168468 174055 168546 174064
rect 168576 174103 168654 174113
rect 168576 174064 168583 174103
rect 168647 174064 168654 174103
rect 168576 173916 168654 174064
rect 169478 174103 169566 174114
rect 169478 174064 169484 174103
rect 169559 174064 169566 174103
rect 169478 174052 169566 174064
rect 168575 173896 168654 173916
rect 169480 173896 169566 174052
rect 168575 173839 168653 173896
rect 168373 173771 168653 173839
rect 166480 173762 166985 173764
rect 168373 173763 168652 173771
rect 167708 173762 168652 173763
rect 166480 173728 168652 173762
rect 166480 173321 168449 173728
rect 168574 173725 168652 173728
rect 166480 173320 167724 173321
rect 166480 170650 166985 173320
rect 167245 173319 167724 173320
rect 169435 170650 169912 173896
rect 170510 172755 171015 174141
rect 189967 174120 190046 174368
rect 193010 174204 193515 174368
rect 192749 174203 193515 174204
rect 190171 174184 193515 174203
rect 190171 174150 190186 174184
rect 192127 174150 193515 174184
rect 190171 174141 193515 174150
rect 190171 174137 192166 174141
rect 189968 174103 190046 174120
rect 189968 174064 189974 174103
rect 190038 174064 190046 174103
rect 189968 174055 190046 174064
rect 190076 174103 190154 174113
rect 190076 174064 190083 174103
rect 190147 174064 190154 174103
rect 192178 174103 192266 174114
rect 192178 174066 192184 174103
rect 190076 173916 190154 174064
rect 190075 173896 190154 173916
rect 192177 174064 192184 174066
rect 192259 174064 192266 174103
rect 190075 173869 190153 173896
rect 189429 173867 190153 173869
rect 188985 173734 190153 173867
rect 192177 173824 192266 174064
rect 192177 173797 192267 173824
rect 188985 172250 189484 173734
rect 190075 173733 190153 173734
rect 192178 173606 192267 173797
rect 192177 173555 192267 173606
rect 192177 173132 192266 173555
rect 192177 173107 192267 173132
rect 192178 172904 192267 173107
rect 188980 170650 189485 172250
rect 192104 170830 192426 172904
rect 193010 172755 193515 174141
rect 169439 170289 169887 170650
rect 192069 170370 192517 170830
rect 168311 151362 168743 151639
rect 168468 151307 168545 151362
rect 168468 151103 168546 151307
rect 170510 151203 171015 151368
rect 189809 151362 190194 151874
rect 168649 151183 171015 151203
rect 168649 151150 168657 151183
rect 168649 151148 168680 151150
rect 169445 151148 171015 151183
rect 168649 151141 171015 151148
rect 168468 151044 168474 151103
rect 168538 151044 168546 151103
rect 168468 151035 168546 151044
rect 168576 151103 168654 151113
rect 168576 151044 168583 151103
rect 168647 151044 168654 151103
rect 168576 150916 168654 151044
rect 169478 151103 169566 151114
rect 169478 151044 169484 151103
rect 169559 151044 169566 151103
rect 169478 151032 169566 151044
rect 168575 150896 168654 150916
rect 169480 150896 169566 151032
rect 168575 150839 168653 150896
rect 168373 150771 168653 150839
rect 166480 150762 166985 150764
rect 168373 150763 168652 150771
rect 167708 150762 168652 150763
rect 166480 150728 168652 150762
rect 166480 150321 168449 150728
rect 168574 150725 168652 150728
rect 166480 150320 167724 150321
rect 166480 147650 166985 150320
rect 167245 150319 167724 150320
rect 169435 147783 169912 150896
rect 170510 149755 171015 151141
rect 189967 151120 190046 151362
rect 193010 151204 193515 151368
rect 192749 151203 193515 151204
rect 190171 151184 193515 151203
rect 190171 151150 190186 151184
rect 192127 151150 193515 151184
rect 190171 151141 193515 151150
rect 190171 151137 192166 151141
rect 189968 151103 190046 151120
rect 189968 151044 189974 151103
rect 190038 151044 190046 151103
rect 189968 151035 190046 151044
rect 190076 151103 190154 151113
rect 190076 151044 190083 151103
rect 190147 151044 190154 151103
rect 192178 151103 192266 151114
rect 192178 151066 192184 151103
rect 190076 150916 190154 151044
rect 190075 150896 190154 150916
rect 192177 151044 192184 151066
rect 192259 151044 192266 151103
rect 190075 150869 190153 150896
rect 189429 150867 190153 150869
rect 188985 150734 190153 150867
rect 192177 150824 192266 151044
rect 192177 150797 192267 150824
rect 188985 149250 189484 150734
rect 190075 150733 190153 150734
rect 192178 150606 192267 150797
rect 192177 150555 192267 150606
rect 192177 150132 192266 150555
rect 192177 150107 192267 150132
rect 192178 149904 192267 150107
rect 169435 147650 169929 147783
rect 188980 147650 189485 149250
rect 192104 148155 192426 149904
rect 193010 149755 193515 151141
rect 169438 147399 169929 147650
rect 192095 147258 192431 148155
rect 168346 128354 168794 128926
rect 168468 128307 168545 128354
rect 168468 128103 168546 128307
rect 170510 128203 171015 128368
rect 189801 128354 190249 128926
rect 168649 128183 171015 128203
rect 168649 128150 168657 128183
rect 168649 128148 168680 128150
rect 169445 128148 171015 128183
rect 168649 128141 171015 128148
rect 168468 128028 168474 128103
rect 168538 128028 168546 128103
rect 168468 128019 168546 128028
rect 168576 128103 168654 128113
rect 168576 128028 168583 128103
rect 168647 128028 168654 128103
rect 168576 127916 168654 128028
rect 169478 128103 169566 128114
rect 169478 128028 169484 128103
rect 169559 128028 169566 128103
rect 169478 128016 169566 128028
rect 168575 127896 168654 127916
rect 169480 127896 169566 128016
rect 168575 127839 168653 127896
rect 168373 127771 168653 127839
rect 166480 127762 166985 127764
rect 168373 127763 168652 127771
rect 167708 127762 168652 127763
rect 166480 127728 168652 127762
rect 166480 127321 168449 127728
rect 168574 127725 168652 127728
rect 166480 127320 167724 127321
rect 166480 124650 166985 127320
rect 167245 127319 167724 127320
rect 169435 124931 169912 127896
rect 170510 126755 171015 128141
rect 189967 128120 190046 128354
rect 193010 128204 193515 128368
rect 192749 128203 193515 128204
rect 190171 128184 193515 128203
rect 190171 128150 190186 128184
rect 192127 128150 193515 128184
rect 190171 128141 193515 128150
rect 190171 128137 192166 128141
rect 189968 128103 190046 128120
rect 189968 128028 189974 128103
rect 190038 128028 190046 128103
rect 189968 128019 190046 128028
rect 190076 128103 190154 128113
rect 190076 128028 190083 128103
rect 190147 128028 190154 128103
rect 192178 128103 192266 128114
rect 192178 128066 192184 128103
rect 190076 127916 190154 128028
rect 190075 127896 190154 127916
rect 192177 128028 192184 128066
rect 192259 128028 192266 128103
rect 190075 127869 190153 127896
rect 189429 127867 190153 127869
rect 188985 127734 190153 127867
rect 192177 127824 192266 128028
rect 192177 127797 192267 127824
rect 188985 126250 189484 127734
rect 190075 127733 190153 127734
rect 192178 127606 192267 127797
rect 192177 127555 192267 127606
rect 192177 127132 192266 127555
rect 192177 127107 192267 127132
rect 192178 126904 192267 127107
rect 169415 124650 169912 124931
rect 188980 124650 189485 126250
rect 192104 124846 192426 126904
rect 193010 126755 193515 128141
rect 169415 124359 169863 124650
rect 192040 124274 192488 124846
rect 168268 105337 168698 105977
rect 168468 105307 168545 105337
rect 168468 105103 168546 105307
rect 170510 105203 171015 105368
rect 189711 105346 190141 105986
rect 168649 105183 171015 105203
rect 168649 105150 168657 105183
rect 168649 105148 168680 105150
rect 169445 105148 171015 105183
rect 168649 105141 171015 105148
rect 168468 104963 168474 105103
rect 168538 104963 168546 105103
rect 168468 104954 168546 104963
rect 168576 105103 168654 105113
rect 168576 104963 168583 105103
rect 168647 104963 168654 105103
rect 168576 104916 168654 104963
rect 169478 105103 169566 105114
rect 169478 104963 169484 105103
rect 169559 104963 169566 105103
rect 169478 104951 169566 104963
rect 168575 104896 168654 104916
rect 169480 104896 169566 104951
rect 168575 104839 168653 104896
rect 168373 104771 168653 104839
rect 166480 104762 166985 104764
rect 168373 104763 168652 104771
rect 167708 104762 168652 104763
rect 166480 104728 168652 104762
rect 166480 104321 168449 104728
rect 168574 104725 168652 104728
rect 166480 104320 167724 104321
rect 166480 101650 166985 104320
rect 167245 104319 167724 104320
rect 169435 101904 169912 104896
rect 170510 103755 171015 105141
rect 189967 105120 190046 105346
rect 193010 105204 193515 105368
rect 192749 105203 193515 105204
rect 190171 105184 193515 105203
rect 190171 105150 190186 105184
rect 192127 105150 193515 105184
rect 190171 105141 193515 105150
rect 190171 105137 192166 105141
rect 189968 105103 190046 105120
rect 189968 104963 189974 105103
rect 190038 104963 190046 105103
rect 189968 104954 190046 104963
rect 190076 105103 190154 105113
rect 190076 104963 190083 105103
rect 190147 104963 190154 105103
rect 192178 105103 192266 105114
rect 192178 105066 192184 105103
rect 190076 104916 190154 104963
rect 190075 104896 190154 104916
rect 192177 104963 192184 105066
rect 192259 104963 192266 105103
rect 190075 104869 190153 104896
rect 189429 104867 190153 104869
rect 188985 104734 190153 104867
rect 192177 104824 192266 104963
rect 192177 104797 192267 104824
rect 188985 103250 189484 104734
rect 190075 104733 190153 104734
rect 192178 104606 192267 104797
rect 192177 104555 192267 104606
rect 192177 104132 192266 104555
rect 192177 104107 192267 104132
rect 192178 103904 192267 104107
rect 169430 101650 169912 101904
rect 188980 101650 189485 103250
rect 192104 102021 192426 103904
rect 193010 103755 193515 105141
rect 192104 101650 192537 102021
rect 169430 101264 169860 101650
rect 192107 101381 192537 101650
rect 168327 82344 168767 82899
rect 189752 82882 190192 82943
rect 189744 82388 190192 82882
rect 168468 82307 168545 82344
rect 168468 82103 168546 82307
rect 170510 82203 171015 82368
rect 189744 82327 190184 82388
rect 168649 82183 171015 82203
rect 168649 82150 168657 82183
rect 168649 82148 168680 82150
rect 169445 82148 171015 82183
rect 168649 82141 171015 82148
rect 168468 81839 168474 82103
rect 168373 81828 168474 81839
rect 168538 81839 168546 82103
rect 168576 82103 168654 82113
rect 168576 81916 168583 82103
rect 168575 81839 168583 81916
rect 168538 81828 168583 81839
rect 168647 81828 168654 82103
rect 169478 82103 169566 82114
rect 169478 81896 169484 82103
rect 168373 81816 168654 81828
rect 169435 81828 169484 81896
rect 169559 81896 169566 82103
rect 169559 81828 169912 81896
rect 168373 81771 168653 81816
rect 166480 81762 166985 81764
rect 168373 81763 168652 81771
rect 167708 81762 168652 81763
rect 166480 81728 168652 81762
rect 166480 81321 168449 81728
rect 168574 81725 168652 81728
rect 166480 81320 167724 81321
rect 166480 78650 166985 81320
rect 167245 81319 167724 81320
rect 169435 78845 169912 81828
rect 170510 80755 171015 82141
rect 189967 82120 190046 82327
rect 193010 82204 193515 82368
rect 192749 82203 193515 82204
rect 190171 82184 193515 82203
rect 190171 82150 190186 82184
rect 192127 82150 193515 82184
rect 190171 82141 193515 82150
rect 190171 82137 192166 82141
rect 189968 82103 190046 82120
rect 189968 81869 189974 82103
rect 189429 81867 189974 81869
rect 188985 81828 189974 81867
rect 190038 81869 190046 82103
rect 190076 82103 190154 82113
rect 190076 81916 190083 82103
rect 190075 81869 190083 81916
rect 190038 81828 190083 81869
rect 190147 81828 190154 82103
rect 192178 82103 192266 82114
rect 192178 82066 192184 82103
rect 188985 81816 190154 81828
rect 192177 81828 192184 82066
rect 192259 81828 192266 82103
rect 192177 81824 192266 81828
rect 188985 81734 190153 81816
rect 192177 81797 192267 81824
rect 188985 80250 189484 81734
rect 190075 81733 190153 81734
rect 192178 81606 192267 81797
rect 192177 81555 192267 81606
rect 192177 81132 192266 81555
rect 192177 81107 192267 81132
rect 192178 80904 192267 81107
rect 169429 78650 169912 78845
rect 188980 78650 189485 80250
rect 192104 78995 192426 80904
rect 193010 80755 193515 82141
rect 169429 78290 169869 78650
rect 192044 78440 192484 78995
rect 168139 59340 168843 60096
rect 168468 59307 168545 59340
rect 168468 59103 168546 59307
rect 170510 59203 171015 59368
rect 189786 59355 191202 59651
rect 168649 59183 171015 59203
rect 168649 59150 168657 59183
rect 168649 59148 168680 59150
rect 169445 59148 171015 59183
rect 168649 59141 171015 59148
rect 166480 58762 166985 58764
rect 167708 58762 168091 58763
rect 166480 58569 168091 58762
rect 168468 58628 168474 59103
rect 168538 58628 168546 59103
rect 168576 59103 168654 59113
rect 168576 58916 168583 59103
rect 168575 58725 168583 58916
rect 168468 58619 168546 58628
rect 168576 58628 168583 58725
rect 168647 58628 168654 59103
rect 169478 59103 169566 59114
rect 169478 58896 169484 59103
rect 168576 58569 168654 58628
rect 166480 58339 168654 58569
rect 169435 58628 169484 58896
rect 169559 58896 169566 59103
rect 169559 58628 169912 58896
rect 166480 58321 168649 58339
rect 166480 58320 167724 58321
rect 168066 58320 168649 58321
rect 166480 55650 166985 58320
rect 167245 58319 167724 58320
rect 169435 55978 169912 58628
rect 170510 57755 171015 59141
rect 189967 59120 190046 59355
rect 193010 59204 193515 59368
rect 192749 59203 193515 59204
rect 190171 59184 193515 59203
rect 190171 59150 190186 59184
rect 192127 59150 193515 59184
rect 190171 59141 193515 59150
rect 190171 59137 192166 59141
rect 189968 59103 190046 59120
rect 189968 58628 189974 59103
rect 190038 58628 190046 59103
rect 190076 59103 190154 59113
rect 190076 58916 190083 59103
rect 189968 58619 190046 58628
rect 190075 58628 190083 58916
rect 190147 58628 190154 59103
rect 192178 59103 192266 59114
rect 192178 59066 192184 59103
rect 192177 58797 192184 59066
rect 190075 58616 190154 58628
rect 192178 58628 192184 58797
rect 192259 58824 192266 59103
rect 192259 58628 192267 58824
rect 190075 58530 190152 58616
rect 192178 58606 192267 58628
rect 188988 58417 190152 58530
rect 188985 58277 190152 58417
rect 192177 58555 192267 58606
rect 188985 58188 190150 58277
rect 188985 57250 189484 58188
rect 192177 58132 192266 58555
rect 192177 58107 192267 58132
rect 192178 57904 192267 58107
rect 169314 55222 170018 55978
rect 188980 55650 189485 57250
rect 192104 55767 192426 57904
rect 193010 57755 193515 59141
rect 192061 55393 192447 55767
rect 167870 36337 168739 36818
rect 168468 36307 168545 36337
rect 168468 36103 168546 36307
rect 170510 36203 171015 36368
rect 189761 36315 190291 36584
rect 168649 36183 171015 36203
rect 168649 36150 168657 36183
rect 168649 36148 168680 36150
rect 169445 36148 171015 36183
rect 168649 36141 171015 36148
rect 168468 35428 168474 36103
rect 168538 35428 168546 36103
rect 168468 35419 168546 35428
rect 168576 36103 168654 36113
rect 168576 35428 168583 36103
rect 168647 35428 168654 36103
rect 168576 35416 168654 35428
rect 169478 36103 169566 36114
rect 169478 35428 169484 36103
rect 169559 35948 169566 36103
rect 169559 35428 169812 35948
rect 169478 35416 169812 35428
rect 170510 35416 171015 36141
rect 189967 36120 190046 36315
rect 193010 36204 193515 36368
rect 192749 36203 193515 36204
rect 190171 36184 193515 36203
rect 190171 36150 190186 36184
rect 192127 36150 193515 36184
rect 190171 36141 193515 36150
rect 190171 36137 192166 36141
rect 189968 36103 190046 36120
rect 189968 35428 189974 36103
rect 190038 35428 190046 36103
rect 189968 35419 190046 35428
rect 190076 36103 190154 36113
rect 190076 35428 190083 36103
rect 190147 35593 190154 36103
rect 192178 36103 192266 36114
rect 190147 35428 190159 35593
rect 190076 35416 190159 35428
rect 192178 35428 192184 36103
rect 192259 35973 192266 36103
rect 192259 35428 192426 35973
rect 192178 35416 192426 35428
rect 193010 35416 193515 36141
rect 166480 34728 166985 34732
rect 168576 34728 168646 35416
rect 169498 34732 169812 35416
rect 190078 35006 190159 35416
rect 166446 34191 168647 34728
rect 166480 32650 166985 34191
rect 169435 33007 169912 34732
rect 188979 34345 190161 35006
rect 192203 34732 192426 35416
rect 188985 34250 189484 34345
rect 169396 32650 169912 33007
rect 188980 32650 189485 34250
rect 192104 32917 192426 34732
rect 169396 32166 169905 32650
rect 192088 32126 192441 32917
rect 167914 13359 168718 13880
rect 168468 13307 168545 13359
rect 168468 13103 168546 13307
rect 170510 13203 171015 13368
rect 189802 13361 190873 13959
rect 168649 13183 171015 13203
rect 168649 13150 168657 13183
rect 168649 13148 168680 13150
rect 169445 13148 171015 13183
rect 168649 13141 171015 13148
rect 166453 3038 167005 10655
rect 168468 3128 168474 13103
rect 168538 3128 168546 13103
rect 168468 3119 168546 3128
rect 168576 13103 168654 13113
rect 168576 3128 168583 13103
rect 168647 3128 168654 13103
rect 168576 3038 168654 3128
rect 169478 13103 169566 13114
rect 169478 3128 169484 13103
rect 169559 3128 169566 13103
rect 170510 12469 171015 13141
rect 189967 13120 190046 13361
rect 193010 13204 193515 13368
rect 192749 13203 193515 13204
rect 190171 13184 193515 13203
rect 190171 13150 190186 13184
rect 192127 13150 193515 13184
rect 190171 13141 193515 13150
rect 190171 13137 192166 13141
rect 189968 13103 190046 13120
rect 169478 3116 169566 3128
rect 166453 2950 168654 3038
rect 188939 3044 189507 10879
rect 189968 3128 189974 13103
rect 190038 3128 190046 13103
rect 189968 3119 190046 3128
rect 190076 13103 190154 13113
rect 190076 3128 190083 13103
rect 190147 3128 190154 13103
rect 190076 3116 190154 3128
rect 192178 13103 192266 13114
rect 192178 3128 192184 13103
rect 192259 3128 192266 13103
rect 192178 3116 192266 3128
rect 193010 3116 193515 13141
rect 190077 3044 190154 3116
rect 166453 2812 168652 2950
rect 188939 2897 190154 3044
rect 188939 2678 190152 2897
use BarePadArray  BarePadArray_0
timestamp 1663654425
transform 1 0 160565 0 1 220400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_1
timestamp 1663654425
transform 1 0 183065 0 1 220400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_2
timestamp 1663654425
transform 1 0 183065 0 1 197400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_3
timestamp 1663654425
transform 1 0 160565 0 1 197400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_4
timestamp 1663654425
transform 1 0 183065 0 1 174400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_5
timestamp 1663654425
transform 1 0 160565 0 1 174400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_6
timestamp 1663654425
transform 1 0 183065 0 1 151400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_7
timestamp 1663654425
transform 1 0 160565 0 1 151400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_8
timestamp 1663654425
transform 1 0 183065 0 1 128400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_9
timestamp 1663654425
transform 1 0 160565 0 1 128400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_10
timestamp 1663654425
transform 1 0 183065 0 1 105400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_11
timestamp 1663654425
transform 1 0 160565 0 1 105400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_12
timestamp 1663654425
transform 1 0 183065 0 1 82400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_13
timestamp 1663654425
transform 1 0 160565 0 1 82400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_14
timestamp 1663654425
transform 1 0 183065 0 1 59400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_15
timestamp 1663654425
transform 1 0 160565 0 1 59400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_16
timestamp 1663654425
transform 1 0 183065 0 1 36400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_17
timestamp 1663654425
transform 1 0 160565 0 1 36400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_18
timestamp 1663654425
transform 1 0 183065 0 1 13400
box -3080 -13385 19420 9615
use BarePadArray  BarePadArray_19
timestamp 1663654425
transform 1 0 160565 0 1 13400
box -3080 -13385 19420 9615
<< end >>
