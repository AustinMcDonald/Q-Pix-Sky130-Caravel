magic
tech sky130B
magscale 1 2
timestamp 1606718285
<< error_p >>
rect -1445 71 -1387 77
rect -1327 71 -1269 77
rect -1209 71 -1151 77
rect -1091 71 -1033 77
rect -973 71 -915 77
rect -855 71 -797 77
rect -737 71 -679 77
rect -619 71 -561 77
rect -501 71 -443 77
rect -383 71 -325 77
rect -265 71 -207 77
rect -147 71 -89 77
rect -29 71 29 77
rect 89 71 147 77
rect 207 71 265 77
rect 325 71 383 77
rect 443 71 501 77
rect 561 71 619 77
rect 679 71 737 77
rect 797 71 855 77
rect 915 71 973 77
rect 1033 71 1091 77
rect 1151 71 1209 77
rect 1269 71 1327 77
rect 1387 71 1445 77
rect -1445 37 -1433 71
rect -1327 37 -1315 71
rect -1209 37 -1197 71
rect -1091 37 -1079 71
rect -973 37 -961 71
rect -855 37 -843 71
rect -737 37 -725 71
rect -619 37 -607 71
rect -501 37 -489 71
rect -383 37 -371 71
rect -265 37 -253 71
rect -147 37 -135 71
rect -29 37 -17 71
rect 89 37 101 71
rect 207 37 219 71
rect 325 37 337 71
rect 443 37 455 71
rect 561 37 573 71
rect 679 37 691 71
rect 797 37 809 71
rect 915 37 927 71
rect 1033 37 1045 71
rect 1151 37 1163 71
rect 1269 37 1281 71
rect 1387 37 1399 71
rect -1445 31 -1387 37
rect -1327 31 -1269 37
rect -1209 31 -1151 37
rect -1091 31 -1033 37
rect -973 31 -915 37
rect -855 31 -797 37
rect -737 31 -679 37
rect -619 31 -561 37
rect -501 31 -443 37
rect -383 31 -325 37
rect -265 31 -207 37
rect -147 31 -89 37
rect -29 31 29 37
rect 89 31 147 37
rect 207 31 265 37
rect 325 31 383 37
rect 443 31 501 37
rect 561 31 619 37
rect 679 31 737 37
rect 797 31 855 37
rect 915 31 973 37
rect 1033 31 1091 37
rect 1151 31 1209 37
rect 1269 31 1327 37
rect 1387 31 1445 37
rect -1445 -37 -1387 -31
rect -1327 -37 -1269 -31
rect -1209 -37 -1151 -31
rect -1091 -37 -1033 -31
rect -973 -37 -915 -31
rect -855 -37 -797 -31
rect -737 -37 -679 -31
rect -619 -37 -561 -31
rect -501 -37 -443 -31
rect -383 -37 -325 -31
rect -265 -37 -207 -31
rect -147 -37 -89 -31
rect -29 -37 29 -31
rect 89 -37 147 -31
rect 207 -37 265 -31
rect 325 -37 383 -31
rect 443 -37 501 -31
rect 561 -37 619 -31
rect 679 -37 737 -31
rect 797 -37 855 -31
rect 915 -37 973 -31
rect 1033 -37 1091 -31
rect 1151 -37 1209 -31
rect 1269 -37 1327 -31
rect 1387 -37 1445 -31
rect -1445 -71 -1433 -37
rect -1327 -71 -1315 -37
rect -1209 -71 -1197 -37
rect -1091 -71 -1079 -37
rect -973 -71 -961 -37
rect -855 -71 -843 -37
rect -737 -71 -725 -37
rect -619 -71 -607 -37
rect -501 -71 -489 -37
rect -383 -71 -371 -37
rect -265 -71 -253 -37
rect -147 -71 -135 -37
rect -29 -71 -17 -37
rect 89 -71 101 -37
rect 207 -71 219 -37
rect 325 -71 337 -37
rect 443 -71 455 -37
rect 561 -71 573 -37
rect 679 -71 691 -37
rect 797 -71 809 -37
rect 915 -71 927 -37
rect 1033 -71 1045 -37
rect 1151 -71 1163 -37
rect 1269 -71 1281 -37
rect 1387 -71 1399 -37
rect -1445 -77 -1387 -71
rect -1327 -77 -1269 -71
rect -1209 -77 -1151 -71
rect -1091 -77 -1033 -71
rect -973 -77 -915 -71
rect -855 -77 -797 -71
rect -737 -77 -679 -71
rect -619 -77 -561 -71
rect -501 -77 -443 -71
rect -383 -77 -325 -71
rect -265 -77 -207 -71
rect -147 -77 -89 -71
rect -29 -77 29 -71
rect 89 -77 147 -71
rect 207 -77 265 -71
rect 325 -77 383 -71
rect 443 -77 501 -71
rect 561 -77 619 -71
rect 679 -77 737 -71
rect 797 -77 855 -71
rect 915 -77 973 -71
rect 1033 -77 1091 -71
rect 1151 -77 1209 -71
rect 1269 -77 1327 -71
rect 1387 -77 1445 -71
<< nwell >>
rect -1642 -937 1642 937
<< pmos >>
rect -1446 118 -1386 718
rect -1328 118 -1268 718
rect -1210 118 -1150 718
rect -1092 118 -1032 718
rect -974 118 -914 718
rect -856 118 -796 718
rect -738 118 -678 718
rect -620 118 -560 718
rect -502 118 -442 718
rect -384 118 -324 718
rect -266 118 -206 718
rect -148 118 -88 718
rect -30 118 30 718
rect 88 118 148 718
rect 206 118 266 718
rect 324 118 384 718
rect 442 118 502 718
rect 560 118 620 718
rect 678 118 738 718
rect 796 118 856 718
rect 914 118 974 718
rect 1032 118 1092 718
rect 1150 118 1210 718
rect 1268 118 1328 718
rect 1386 118 1446 718
rect -1446 -718 -1386 -118
rect -1328 -718 -1268 -118
rect -1210 -718 -1150 -118
rect -1092 -718 -1032 -118
rect -974 -718 -914 -118
rect -856 -718 -796 -118
rect -738 -718 -678 -118
rect -620 -718 -560 -118
rect -502 -718 -442 -118
rect -384 -718 -324 -118
rect -266 -718 -206 -118
rect -148 -718 -88 -118
rect -30 -718 30 -118
rect 88 -718 148 -118
rect 206 -718 266 -118
rect 324 -718 384 -118
rect 442 -718 502 -118
rect 560 -718 620 -118
rect 678 -718 738 -118
rect 796 -718 856 -118
rect 914 -718 974 -118
rect 1032 -718 1092 -118
rect 1150 -718 1210 -118
rect 1268 -718 1328 -118
rect 1386 -718 1446 -118
<< pdiff >>
rect -1504 706 -1446 718
rect -1504 130 -1492 706
rect -1458 130 -1446 706
rect -1504 118 -1446 130
rect -1386 706 -1328 718
rect -1386 130 -1374 706
rect -1340 130 -1328 706
rect -1386 118 -1328 130
rect -1268 706 -1210 718
rect -1268 130 -1256 706
rect -1222 130 -1210 706
rect -1268 118 -1210 130
rect -1150 706 -1092 718
rect -1150 130 -1138 706
rect -1104 130 -1092 706
rect -1150 118 -1092 130
rect -1032 706 -974 718
rect -1032 130 -1020 706
rect -986 130 -974 706
rect -1032 118 -974 130
rect -914 706 -856 718
rect -914 130 -902 706
rect -868 130 -856 706
rect -914 118 -856 130
rect -796 706 -738 718
rect -796 130 -784 706
rect -750 130 -738 706
rect -796 118 -738 130
rect -678 706 -620 718
rect -678 130 -666 706
rect -632 130 -620 706
rect -678 118 -620 130
rect -560 706 -502 718
rect -560 130 -548 706
rect -514 130 -502 706
rect -560 118 -502 130
rect -442 706 -384 718
rect -442 130 -430 706
rect -396 130 -384 706
rect -442 118 -384 130
rect -324 706 -266 718
rect -324 130 -312 706
rect -278 130 -266 706
rect -324 118 -266 130
rect -206 706 -148 718
rect -206 130 -194 706
rect -160 130 -148 706
rect -206 118 -148 130
rect -88 706 -30 718
rect -88 130 -76 706
rect -42 130 -30 706
rect -88 118 -30 130
rect 30 706 88 718
rect 30 130 42 706
rect 76 130 88 706
rect 30 118 88 130
rect 148 706 206 718
rect 148 130 160 706
rect 194 130 206 706
rect 148 118 206 130
rect 266 706 324 718
rect 266 130 278 706
rect 312 130 324 706
rect 266 118 324 130
rect 384 706 442 718
rect 384 130 396 706
rect 430 130 442 706
rect 384 118 442 130
rect 502 706 560 718
rect 502 130 514 706
rect 548 130 560 706
rect 502 118 560 130
rect 620 706 678 718
rect 620 130 632 706
rect 666 130 678 706
rect 620 118 678 130
rect 738 706 796 718
rect 738 130 750 706
rect 784 130 796 706
rect 738 118 796 130
rect 856 706 914 718
rect 856 130 868 706
rect 902 130 914 706
rect 856 118 914 130
rect 974 706 1032 718
rect 974 130 986 706
rect 1020 130 1032 706
rect 974 118 1032 130
rect 1092 706 1150 718
rect 1092 130 1104 706
rect 1138 130 1150 706
rect 1092 118 1150 130
rect 1210 706 1268 718
rect 1210 130 1222 706
rect 1256 130 1268 706
rect 1210 118 1268 130
rect 1328 706 1386 718
rect 1328 130 1340 706
rect 1374 130 1386 706
rect 1328 118 1386 130
rect 1446 706 1504 718
rect 1446 130 1458 706
rect 1492 130 1504 706
rect 1446 118 1504 130
rect -1504 -130 -1446 -118
rect -1504 -706 -1492 -130
rect -1458 -706 -1446 -130
rect -1504 -718 -1446 -706
rect -1386 -130 -1328 -118
rect -1386 -706 -1374 -130
rect -1340 -706 -1328 -130
rect -1386 -718 -1328 -706
rect -1268 -130 -1210 -118
rect -1268 -706 -1256 -130
rect -1222 -706 -1210 -130
rect -1268 -718 -1210 -706
rect -1150 -130 -1092 -118
rect -1150 -706 -1138 -130
rect -1104 -706 -1092 -130
rect -1150 -718 -1092 -706
rect -1032 -130 -974 -118
rect -1032 -706 -1020 -130
rect -986 -706 -974 -130
rect -1032 -718 -974 -706
rect -914 -130 -856 -118
rect -914 -706 -902 -130
rect -868 -706 -856 -130
rect -914 -718 -856 -706
rect -796 -130 -738 -118
rect -796 -706 -784 -130
rect -750 -706 -738 -130
rect -796 -718 -738 -706
rect -678 -130 -620 -118
rect -678 -706 -666 -130
rect -632 -706 -620 -130
rect -678 -718 -620 -706
rect -560 -130 -502 -118
rect -560 -706 -548 -130
rect -514 -706 -502 -130
rect -560 -718 -502 -706
rect -442 -130 -384 -118
rect -442 -706 -430 -130
rect -396 -706 -384 -130
rect -442 -718 -384 -706
rect -324 -130 -266 -118
rect -324 -706 -312 -130
rect -278 -706 -266 -130
rect -324 -718 -266 -706
rect -206 -130 -148 -118
rect -206 -706 -194 -130
rect -160 -706 -148 -130
rect -206 -718 -148 -706
rect -88 -130 -30 -118
rect -88 -706 -76 -130
rect -42 -706 -30 -130
rect -88 -718 -30 -706
rect 30 -130 88 -118
rect 30 -706 42 -130
rect 76 -706 88 -130
rect 30 -718 88 -706
rect 148 -130 206 -118
rect 148 -706 160 -130
rect 194 -706 206 -130
rect 148 -718 206 -706
rect 266 -130 324 -118
rect 266 -706 278 -130
rect 312 -706 324 -130
rect 266 -718 324 -706
rect 384 -130 442 -118
rect 384 -706 396 -130
rect 430 -706 442 -130
rect 384 -718 442 -706
rect 502 -130 560 -118
rect 502 -706 514 -130
rect 548 -706 560 -130
rect 502 -718 560 -706
rect 620 -130 678 -118
rect 620 -706 632 -130
rect 666 -706 678 -130
rect 620 -718 678 -706
rect 738 -130 796 -118
rect 738 -706 750 -130
rect 784 -706 796 -130
rect 738 -718 796 -706
rect 856 -130 914 -118
rect 856 -706 868 -130
rect 902 -706 914 -130
rect 856 -718 914 -706
rect 974 -130 1032 -118
rect 974 -706 986 -130
rect 1020 -706 1032 -130
rect 974 -718 1032 -706
rect 1092 -130 1150 -118
rect 1092 -706 1104 -130
rect 1138 -706 1150 -130
rect 1092 -718 1150 -706
rect 1210 -130 1268 -118
rect 1210 -706 1222 -130
rect 1256 -706 1268 -130
rect 1210 -718 1268 -706
rect 1328 -130 1386 -118
rect 1328 -706 1340 -130
rect 1374 -706 1386 -130
rect 1328 -718 1386 -706
rect 1446 -130 1504 -118
rect 1446 -706 1458 -130
rect 1492 -706 1504 -130
rect 1446 -718 1504 -706
<< pdiffc >>
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect -1492 -706 -1458 -130
rect -1374 -706 -1340 -130
rect -1256 -706 -1222 -130
rect -1138 -706 -1104 -130
rect -1020 -706 -986 -130
rect -902 -706 -868 -130
rect -784 -706 -750 -130
rect -666 -706 -632 -130
rect -548 -706 -514 -130
rect -430 -706 -396 -130
rect -312 -706 -278 -130
rect -194 -706 -160 -130
rect -76 -706 -42 -130
rect 42 -706 76 -130
rect 160 -706 194 -130
rect 278 -706 312 -130
rect 396 -706 430 -130
rect 514 -706 548 -130
rect 632 -706 666 -130
rect 750 -706 784 -130
rect 868 -706 902 -130
rect 986 -706 1020 -130
rect 1104 -706 1138 -130
rect 1222 -706 1256 -130
rect 1340 -706 1374 -130
rect 1458 -706 1492 -130
<< nsubdiff >>
rect -1606 867 -1510 901
rect 1510 867 1606 901
rect -1606 805 -1572 867
rect 1572 805 1606 867
rect -1606 -867 -1572 -805
rect 1572 -867 1606 -805
rect -1606 -901 -1510 -867
rect 1510 -901 1606 -867
<< nsubdiffcont >>
rect -1510 867 1510 901
rect -1606 -805 -1572 805
rect 1572 -805 1606 805
rect -1510 -901 1510 -867
<< poly >>
rect -1449 749 -1383 815
rect -1331 749 -1265 815
rect -1213 749 -1147 815
rect -1095 749 -1029 815
rect -977 749 -911 815
rect -859 749 -793 815
rect -741 749 -675 815
rect -623 749 -557 815
rect -505 749 -439 815
rect -387 749 -321 815
rect -269 749 -203 815
rect -151 749 -85 815
rect -33 749 33 815
rect 85 749 151 815
rect 203 749 269 815
rect 321 749 387 815
rect 439 749 505 815
rect 557 749 623 815
rect 675 749 741 815
rect 793 749 859 815
rect 911 749 977 815
rect 1029 749 1095 815
rect 1147 749 1213 815
rect 1265 749 1331 815
rect 1383 749 1449 815
rect -1446 718 -1386 749
rect -1328 718 -1268 749
rect -1210 718 -1150 749
rect -1092 718 -1032 749
rect -974 718 -914 749
rect -856 718 -796 749
rect -738 718 -678 749
rect -620 718 -560 749
rect -502 718 -442 749
rect -384 718 -324 749
rect -266 718 -206 749
rect -148 718 -88 749
rect -30 718 30 749
rect 88 718 148 749
rect 206 718 266 749
rect 324 718 384 749
rect 442 718 502 749
rect 560 718 620 749
rect 678 718 738 749
rect 796 718 856 749
rect 914 718 974 749
rect 1032 718 1092 749
rect 1150 718 1210 749
rect 1268 718 1328 749
rect 1386 718 1446 749
rect -1446 87 -1386 118
rect -1328 87 -1268 118
rect -1210 87 -1150 118
rect -1092 87 -1032 118
rect -974 87 -914 118
rect -856 87 -796 118
rect -738 87 -678 118
rect -620 87 -560 118
rect -502 87 -442 118
rect -384 87 -324 118
rect -266 87 -206 118
rect -148 87 -88 118
rect -30 87 30 118
rect 88 87 148 118
rect 206 87 266 118
rect 324 87 384 118
rect 442 87 502 118
rect 560 87 620 118
rect 678 87 738 118
rect 796 87 856 118
rect 914 87 974 118
rect 1032 87 1092 118
rect 1150 87 1210 118
rect 1268 87 1328 118
rect 1386 87 1446 118
rect -1449 71 -1383 87
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1449 21 -1383 37
rect -1331 71 -1265 87
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1331 21 -1265 37
rect -1213 71 -1147 87
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1213 21 -1147 37
rect -1095 71 -1029 87
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -1095 21 -1029 37
rect -977 71 -911 87
rect -977 37 -961 71
rect -927 37 -911 71
rect -977 21 -911 37
rect -859 71 -793 87
rect -859 37 -843 71
rect -809 37 -793 71
rect -859 21 -793 37
rect -741 71 -675 87
rect -741 37 -725 71
rect -691 37 -675 71
rect -741 21 -675 37
rect -623 71 -557 87
rect -623 37 -607 71
rect -573 37 -557 71
rect -623 21 -557 37
rect -505 71 -439 87
rect -505 37 -489 71
rect -455 37 -439 71
rect -505 21 -439 37
rect -387 71 -321 87
rect -387 37 -371 71
rect -337 37 -321 71
rect -387 21 -321 37
rect -269 71 -203 87
rect -269 37 -253 71
rect -219 37 -203 71
rect -269 21 -203 37
rect -151 71 -85 87
rect -151 37 -135 71
rect -101 37 -85 71
rect -151 21 -85 37
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect 85 71 151 87
rect 85 37 101 71
rect 135 37 151 71
rect 85 21 151 37
rect 203 71 269 87
rect 203 37 219 71
rect 253 37 269 71
rect 203 21 269 37
rect 321 71 387 87
rect 321 37 337 71
rect 371 37 387 71
rect 321 21 387 37
rect 439 71 505 87
rect 439 37 455 71
rect 489 37 505 71
rect 439 21 505 37
rect 557 71 623 87
rect 557 37 573 71
rect 607 37 623 71
rect 557 21 623 37
rect 675 71 741 87
rect 675 37 691 71
rect 725 37 741 71
rect 675 21 741 37
rect 793 71 859 87
rect 793 37 809 71
rect 843 37 859 71
rect 793 21 859 37
rect 911 71 977 87
rect 911 37 927 71
rect 961 37 977 71
rect 911 21 977 37
rect 1029 71 1095 87
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1029 21 1095 37
rect 1147 71 1213 87
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1147 21 1213 37
rect 1265 71 1331 87
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1265 21 1331 37
rect 1383 71 1449 87
rect 1383 37 1399 71
rect 1433 37 1449 71
rect 1383 21 1449 37
rect -1449 -37 -1383 -21
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1449 -87 -1383 -71
rect -1331 -37 -1265 -21
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1331 -87 -1265 -71
rect -1213 -37 -1147 -21
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1213 -87 -1147 -71
rect -1095 -37 -1029 -21
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -1095 -87 -1029 -71
rect -977 -37 -911 -21
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -977 -87 -911 -71
rect -859 -37 -793 -21
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -859 -87 -793 -71
rect -741 -37 -675 -21
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -741 -87 -675 -71
rect -623 -37 -557 -21
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -623 -87 -557 -71
rect -505 -37 -439 -21
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -505 -87 -439 -71
rect -387 -37 -321 -21
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -387 -87 -321 -71
rect -269 -37 -203 -21
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -269 -87 -203 -71
rect -151 -37 -85 -21
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -151 -87 -85 -71
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect 85 -37 151 -21
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 85 -87 151 -71
rect 203 -37 269 -21
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 203 -87 269 -71
rect 321 -37 387 -21
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 321 -87 387 -71
rect 439 -37 505 -21
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 439 -87 505 -71
rect 557 -37 623 -21
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 557 -87 623 -71
rect 675 -37 741 -21
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 675 -87 741 -71
rect 793 -37 859 -21
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 793 -87 859 -71
rect 911 -37 977 -21
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 911 -87 977 -71
rect 1029 -37 1095 -21
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1029 -87 1095 -71
rect 1147 -37 1213 -21
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1147 -87 1213 -71
rect 1265 -37 1331 -21
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1265 -87 1331 -71
rect 1383 -37 1449 -21
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect 1383 -87 1449 -71
rect -1446 -118 -1386 -87
rect -1328 -118 -1268 -87
rect -1210 -118 -1150 -87
rect -1092 -118 -1032 -87
rect -974 -118 -914 -87
rect -856 -118 -796 -87
rect -738 -118 -678 -87
rect -620 -118 -560 -87
rect -502 -118 -442 -87
rect -384 -118 -324 -87
rect -266 -118 -206 -87
rect -148 -118 -88 -87
rect -30 -118 30 -87
rect 88 -118 148 -87
rect 206 -118 266 -87
rect 324 -118 384 -87
rect 442 -118 502 -87
rect 560 -118 620 -87
rect 678 -118 738 -87
rect 796 -118 856 -87
rect 914 -118 974 -87
rect 1032 -118 1092 -87
rect 1150 -118 1210 -87
rect 1268 -118 1328 -87
rect 1386 -118 1446 -87
rect -1446 -749 -1386 -718
rect -1328 -749 -1268 -718
rect -1210 -749 -1150 -718
rect -1092 -749 -1032 -718
rect -974 -749 -914 -718
rect -856 -749 -796 -718
rect -738 -749 -678 -718
rect -620 -749 -560 -718
rect -502 -749 -442 -718
rect -384 -749 -324 -718
rect -266 -749 -206 -718
rect -148 -749 -88 -718
rect -30 -749 30 -718
rect 88 -749 148 -718
rect 206 -749 266 -718
rect 324 -749 384 -718
rect 442 -749 502 -718
rect 560 -749 620 -718
rect 678 -749 738 -718
rect 796 -749 856 -718
rect 914 -749 974 -718
rect 1032 -749 1092 -718
rect 1150 -749 1210 -718
rect 1268 -749 1328 -718
rect 1386 -749 1446 -718
rect -1449 -815 -1383 -749
rect -1331 -815 -1265 -749
rect -1213 -815 -1147 -749
rect -1095 -815 -1029 -749
rect -977 -815 -911 -749
rect -859 -815 -793 -749
rect -741 -815 -675 -749
rect -623 -815 -557 -749
rect -505 -815 -439 -749
rect -387 -815 -321 -749
rect -269 -815 -203 -749
rect -151 -815 -85 -749
rect -33 -815 33 -749
rect 85 -815 151 -749
rect 203 -815 269 -749
rect 321 -815 387 -749
rect 439 -815 505 -749
rect 557 -815 623 -749
rect 675 -815 741 -749
rect 793 -815 859 -749
rect 911 -815 977 -749
rect 1029 -815 1095 -749
rect 1147 -815 1213 -749
rect 1265 -815 1331 -749
rect 1383 -815 1449 -749
<< polycont >>
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
<< locali >>
rect -1606 867 -1510 901
rect 1510 867 1606 901
rect -1606 805 -1572 867
rect 1572 805 1606 867
rect -1492 706 -1458 722
rect -1492 114 -1458 130
rect -1374 706 -1340 722
rect -1374 114 -1340 130
rect -1256 706 -1222 722
rect -1256 114 -1222 130
rect -1138 706 -1104 722
rect -1138 114 -1104 130
rect -1020 706 -986 722
rect -1020 114 -986 130
rect -902 706 -868 722
rect -902 114 -868 130
rect -784 706 -750 722
rect -784 114 -750 130
rect -666 706 -632 722
rect -666 114 -632 130
rect -548 706 -514 722
rect -548 114 -514 130
rect -430 706 -396 722
rect -430 114 -396 130
rect -312 706 -278 722
rect -312 114 -278 130
rect -194 706 -160 722
rect -194 114 -160 130
rect -76 706 -42 722
rect -76 114 -42 130
rect 42 706 76 722
rect 42 114 76 130
rect 160 706 194 722
rect 160 114 194 130
rect 278 706 312 722
rect 278 114 312 130
rect 396 706 430 722
rect 396 114 430 130
rect 514 706 548 722
rect 514 114 548 130
rect 632 706 666 722
rect 632 114 666 130
rect 750 706 784 722
rect 750 114 784 130
rect 868 706 902 722
rect 868 114 902 130
rect 986 706 1020 722
rect 986 114 1020 130
rect 1104 706 1138 722
rect 1104 114 1138 130
rect 1222 706 1256 722
rect 1222 114 1256 130
rect 1340 706 1374 722
rect 1340 114 1374 130
rect 1458 706 1492 722
rect 1458 114 1492 130
rect -1449 37 -1433 71
rect -1399 37 -1383 71
rect -1331 37 -1315 71
rect -1281 37 -1265 71
rect -1213 37 -1197 71
rect -1163 37 -1147 71
rect -1095 37 -1079 71
rect -1045 37 -1029 71
rect -977 37 -961 71
rect -927 37 -911 71
rect -859 37 -843 71
rect -809 37 -793 71
rect -741 37 -725 71
rect -691 37 -675 71
rect -623 37 -607 71
rect -573 37 -557 71
rect -505 37 -489 71
rect -455 37 -439 71
rect -387 37 -371 71
rect -337 37 -321 71
rect -269 37 -253 71
rect -219 37 -203 71
rect -151 37 -135 71
rect -101 37 -85 71
rect -33 37 -17 71
rect 17 37 33 71
rect 85 37 101 71
rect 135 37 151 71
rect 203 37 219 71
rect 253 37 269 71
rect 321 37 337 71
rect 371 37 387 71
rect 439 37 455 71
rect 489 37 505 71
rect 557 37 573 71
rect 607 37 623 71
rect 675 37 691 71
rect 725 37 741 71
rect 793 37 809 71
rect 843 37 859 71
rect 911 37 927 71
rect 961 37 977 71
rect 1029 37 1045 71
rect 1079 37 1095 71
rect 1147 37 1163 71
rect 1197 37 1213 71
rect 1265 37 1281 71
rect 1315 37 1331 71
rect 1383 37 1399 71
rect 1433 37 1449 71
rect -1449 -71 -1433 -37
rect -1399 -71 -1383 -37
rect -1331 -71 -1315 -37
rect -1281 -71 -1265 -37
rect -1213 -71 -1197 -37
rect -1163 -71 -1147 -37
rect -1095 -71 -1079 -37
rect -1045 -71 -1029 -37
rect -977 -71 -961 -37
rect -927 -71 -911 -37
rect -859 -71 -843 -37
rect -809 -71 -793 -37
rect -741 -71 -725 -37
rect -691 -71 -675 -37
rect -623 -71 -607 -37
rect -573 -71 -557 -37
rect -505 -71 -489 -37
rect -455 -71 -439 -37
rect -387 -71 -371 -37
rect -337 -71 -321 -37
rect -269 -71 -253 -37
rect -219 -71 -203 -37
rect -151 -71 -135 -37
rect -101 -71 -85 -37
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect 85 -71 101 -37
rect 135 -71 151 -37
rect 203 -71 219 -37
rect 253 -71 269 -37
rect 321 -71 337 -37
rect 371 -71 387 -37
rect 439 -71 455 -37
rect 489 -71 505 -37
rect 557 -71 573 -37
rect 607 -71 623 -37
rect 675 -71 691 -37
rect 725 -71 741 -37
rect 793 -71 809 -37
rect 843 -71 859 -37
rect 911 -71 927 -37
rect 961 -71 977 -37
rect 1029 -71 1045 -37
rect 1079 -71 1095 -37
rect 1147 -71 1163 -37
rect 1197 -71 1213 -37
rect 1265 -71 1281 -37
rect 1315 -71 1331 -37
rect 1383 -71 1399 -37
rect 1433 -71 1449 -37
rect -1492 -130 -1458 -114
rect -1492 -722 -1458 -706
rect -1374 -130 -1340 -114
rect -1374 -722 -1340 -706
rect -1256 -130 -1222 -114
rect -1256 -722 -1222 -706
rect -1138 -130 -1104 -114
rect -1138 -722 -1104 -706
rect -1020 -130 -986 -114
rect -1020 -722 -986 -706
rect -902 -130 -868 -114
rect -902 -722 -868 -706
rect -784 -130 -750 -114
rect -784 -722 -750 -706
rect -666 -130 -632 -114
rect -666 -722 -632 -706
rect -548 -130 -514 -114
rect -548 -722 -514 -706
rect -430 -130 -396 -114
rect -430 -722 -396 -706
rect -312 -130 -278 -114
rect -312 -722 -278 -706
rect -194 -130 -160 -114
rect -194 -722 -160 -706
rect -76 -130 -42 -114
rect -76 -722 -42 -706
rect 42 -130 76 -114
rect 42 -722 76 -706
rect 160 -130 194 -114
rect 160 -722 194 -706
rect 278 -130 312 -114
rect 278 -722 312 -706
rect 396 -130 430 -114
rect 396 -722 430 -706
rect 514 -130 548 -114
rect 514 -722 548 -706
rect 632 -130 666 -114
rect 632 -722 666 -706
rect 750 -130 784 -114
rect 750 -722 784 -706
rect 868 -130 902 -114
rect 868 -722 902 -706
rect 986 -130 1020 -114
rect 986 -722 1020 -706
rect 1104 -130 1138 -114
rect 1104 -722 1138 -706
rect 1222 -130 1256 -114
rect 1222 -722 1256 -706
rect 1340 -130 1374 -114
rect 1340 -722 1374 -706
rect 1458 -130 1492 -114
rect 1458 -722 1492 -706
rect -1606 -867 -1572 -805
rect 1572 -867 1606 -805
rect -1606 -901 -1510 -867
rect 1510 -901 1606 -867
<< viali >>
rect -1492 130 -1458 706
rect -1374 130 -1340 706
rect -1256 130 -1222 706
rect -1138 130 -1104 706
rect -1020 130 -986 706
rect -902 130 -868 706
rect -784 130 -750 706
rect -666 130 -632 706
rect -548 130 -514 706
rect -430 130 -396 706
rect -312 130 -278 706
rect -194 130 -160 706
rect -76 130 -42 706
rect 42 130 76 706
rect 160 130 194 706
rect 278 130 312 706
rect 396 130 430 706
rect 514 130 548 706
rect 632 130 666 706
rect 750 130 784 706
rect 868 130 902 706
rect 986 130 1020 706
rect 1104 130 1138 706
rect 1222 130 1256 706
rect 1340 130 1374 706
rect 1458 130 1492 706
rect -1433 37 -1399 71
rect -1315 37 -1281 71
rect -1197 37 -1163 71
rect -1079 37 -1045 71
rect -961 37 -927 71
rect -843 37 -809 71
rect -725 37 -691 71
rect -607 37 -573 71
rect -489 37 -455 71
rect -371 37 -337 71
rect -253 37 -219 71
rect -135 37 -101 71
rect -17 37 17 71
rect 101 37 135 71
rect 219 37 253 71
rect 337 37 371 71
rect 455 37 489 71
rect 573 37 607 71
rect 691 37 725 71
rect 809 37 843 71
rect 927 37 961 71
rect 1045 37 1079 71
rect 1163 37 1197 71
rect 1281 37 1315 71
rect 1399 37 1433 71
rect -1433 -71 -1399 -37
rect -1315 -71 -1281 -37
rect -1197 -71 -1163 -37
rect -1079 -71 -1045 -37
rect -961 -71 -927 -37
rect -843 -71 -809 -37
rect -725 -71 -691 -37
rect -607 -71 -573 -37
rect -489 -71 -455 -37
rect -371 -71 -337 -37
rect -253 -71 -219 -37
rect -135 -71 -101 -37
rect -17 -71 17 -37
rect 101 -71 135 -37
rect 219 -71 253 -37
rect 337 -71 371 -37
rect 455 -71 489 -37
rect 573 -71 607 -37
rect 691 -71 725 -37
rect 809 -71 843 -37
rect 927 -71 961 -37
rect 1045 -71 1079 -37
rect 1163 -71 1197 -37
rect 1281 -71 1315 -37
rect 1399 -71 1433 -37
rect -1492 -706 -1458 -130
rect -1374 -706 -1340 -130
rect -1256 -706 -1222 -130
rect -1138 -706 -1104 -130
rect -1020 -706 -986 -130
rect -902 -706 -868 -130
rect -784 -706 -750 -130
rect -666 -706 -632 -130
rect -548 -706 -514 -130
rect -430 -706 -396 -130
rect -312 -706 -278 -130
rect -194 -706 -160 -130
rect -76 -706 -42 -130
rect 42 -706 76 -130
rect 160 -706 194 -130
rect 278 -706 312 -130
rect 396 -706 430 -130
rect 514 -706 548 -130
rect 632 -706 666 -130
rect 750 -706 784 -130
rect 868 -706 902 -130
rect 986 -706 1020 -130
rect 1104 -706 1138 -130
rect 1222 -706 1256 -130
rect 1340 -706 1374 -130
rect 1458 -706 1492 -130
<< metal1 >>
rect -1498 706 -1452 718
rect -1498 130 -1492 706
rect -1458 130 -1452 706
rect -1498 118 -1452 130
rect -1380 706 -1334 718
rect -1380 130 -1374 706
rect -1340 130 -1334 706
rect -1380 118 -1334 130
rect -1262 706 -1216 718
rect -1262 130 -1256 706
rect -1222 130 -1216 706
rect -1262 118 -1216 130
rect -1144 706 -1098 718
rect -1144 130 -1138 706
rect -1104 130 -1098 706
rect -1144 118 -1098 130
rect -1026 706 -980 718
rect -1026 130 -1020 706
rect -986 130 -980 706
rect -1026 118 -980 130
rect -908 706 -862 718
rect -908 130 -902 706
rect -868 130 -862 706
rect -908 118 -862 130
rect -790 706 -744 718
rect -790 130 -784 706
rect -750 130 -744 706
rect -790 118 -744 130
rect -672 706 -626 718
rect -672 130 -666 706
rect -632 130 -626 706
rect -672 118 -626 130
rect -554 706 -508 718
rect -554 130 -548 706
rect -514 130 -508 706
rect -554 118 -508 130
rect -436 706 -390 718
rect -436 130 -430 706
rect -396 130 -390 706
rect -436 118 -390 130
rect -318 706 -272 718
rect -318 130 -312 706
rect -278 130 -272 706
rect -318 118 -272 130
rect -200 706 -154 718
rect -200 130 -194 706
rect -160 130 -154 706
rect -200 118 -154 130
rect -82 706 -36 718
rect -82 130 -76 706
rect -42 130 -36 706
rect -82 118 -36 130
rect 36 706 82 718
rect 36 130 42 706
rect 76 130 82 706
rect 36 118 82 130
rect 154 706 200 718
rect 154 130 160 706
rect 194 130 200 706
rect 154 118 200 130
rect 272 706 318 718
rect 272 130 278 706
rect 312 130 318 706
rect 272 118 318 130
rect 390 706 436 718
rect 390 130 396 706
rect 430 130 436 706
rect 390 118 436 130
rect 508 706 554 718
rect 508 130 514 706
rect 548 130 554 706
rect 508 118 554 130
rect 626 706 672 718
rect 626 130 632 706
rect 666 130 672 706
rect 626 118 672 130
rect 744 706 790 718
rect 744 130 750 706
rect 784 130 790 706
rect 744 118 790 130
rect 862 706 908 718
rect 862 130 868 706
rect 902 130 908 706
rect 862 118 908 130
rect 980 706 1026 718
rect 980 130 986 706
rect 1020 130 1026 706
rect 980 118 1026 130
rect 1098 706 1144 718
rect 1098 130 1104 706
rect 1138 130 1144 706
rect 1098 118 1144 130
rect 1216 706 1262 718
rect 1216 130 1222 706
rect 1256 130 1262 706
rect 1216 118 1262 130
rect 1334 706 1380 718
rect 1334 130 1340 706
rect 1374 130 1380 706
rect 1334 118 1380 130
rect 1452 706 1498 718
rect 1452 130 1458 706
rect 1492 130 1498 706
rect 1452 118 1498 130
rect -1445 71 -1387 77
rect -1445 37 -1433 71
rect -1399 37 -1387 71
rect -1445 31 -1387 37
rect -1327 71 -1269 77
rect -1327 37 -1315 71
rect -1281 37 -1269 71
rect -1327 31 -1269 37
rect -1209 71 -1151 77
rect -1209 37 -1197 71
rect -1163 37 -1151 71
rect -1209 31 -1151 37
rect -1091 71 -1033 77
rect -1091 37 -1079 71
rect -1045 37 -1033 71
rect -1091 31 -1033 37
rect -973 71 -915 77
rect -973 37 -961 71
rect -927 37 -915 71
rect -973 31 -915 37
rect -855 71 -797 77
rect -855 37 -843 71
rect -809 37 -797 71
rect -855 31 -797 37
rect -737 71 -679 77
rect -737 37 -725 71
rect -691 37 -679 71
rect -737 31 -679 37
rect -619 71 -561 77
rect -619 37 -607 71
rect -573 37 -561 71
rect -619 31 -561 37
rect -501 71 -443 77
rect -501 37 -489 71
rect -455 37 -443 71
rect -501 31 -443 37
rect -383 71 -325 77
rect -383 37 -371 71
rect -337 37 -325 71
rect -383 31 -325 37
rect -265 71 -207 77
rect -265 37 -253 71
rect -219 37 -207 71
rect -265 31 -207 37
rect -147 71 -89 77
rect -147 37 -135 71
rect -101 37 -89 71
rect -147 31 -89 37
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect 89 71 147 77
rect 89 37 101 71
rect 135 37 147 71
rect 89 31 147 37
rect 207 71 265 77
rect 207 37 219 71
rect 253 37 265 71
rect 207 31 265 37
rect 325 71 383 77
rect 325 37 337 71
rect 371 37 383 71
rect 325 31 383 37
rect 443 71 501 77
rect 443 37 455 71
rect 489 37 501 71
rect 443 31 501 37
rect 561 71 619 77
rect 561 37 573 71
rect 607 37 619 71
rect 561 31 619 37
rect 679 71 737 77
rect 679 37 691 71
rect 725 37 737 71
rect 679 31 737 37
rect 797 71 855 77
rect 797 37 809 71
rect 843 37 855 71
rect 797 31 855 37
rect 915 71 973 77
rect 915 37 927 71
rect 961 37 973 71
rect 915 31 973 37
rect 1033 71 1091 77
rect 1033 37 1045 71
rect 1079 37 1091 71
rect 1033 31 1091 37
rect 1151 71 1209 77
rect 1151 37 1163 71
rect 1197 37 1209 71
rect 1151 31 1209 37
rect 1269 71 1327 77
rect 1269 37 1281 71
rect 1315 37 1327 71
rect 1269 31 1327 37
rect 1387 71 1445 77
rect 1387 37 1399 71
rect 1433 37 1445 71
rect 1387 31 1445 37
rect -1445 -37 -1387 -31
rect -1445 -71 -1433 -37
rect -1399 -71 -1387 -37
rect -1445 -77 -1387 -71
rect -1327 -37 -1269 -31
rect -1327 -71 -1315 -37
rect -1281 -71 -1269 -37
rect -1327 -77 -1269 -71
rect -1209 -37 -1151 -31
rect -1209 -71 -1197 -37
rect -1163 -71 -1151 -37
rect -1209 -77 -1151 -71
rect -1091 -37 -1033 -31
rect -1091 -71 -1079 -37
rect -1045 -71 -1033 -37
rect -1091 -77 -1033 -71
rect -973 -37 -915 -31
rect -973 -71 -961 -37
rect -927 -71 -915 -37
rect -973 -77 -915 -71
rect -855 -37 -797 -31
rect -855 -71 -843 -37
rect -809 -71 -797 -37
rect -855 -77 -797 -71
rect -737 -37 -679 -31
rect -737 -71 -725 -37
rect -691 -71 -679 -37
rect -737 -77 -679 -71
rect -619 -37 -561 -31
rect -619 -71 -607 -37
rect -573 -71 -561 -37
rect -619 -77 -561 -71
rect -501 -37 -443 -31
rect -501 -71 -489 -37
rect -455 -71 -443 -37
rect -501 -77 -443 -71
rect -383 -37 -325 -31
rect -383 -71 -371 -37
rect -337 -71 -325 -37
rect -383 -77 -325 -71
rect -265 -37 -207 -31
rect -265 -71 -253 -37
rect -219 -71 -207 -37
rect -265 -77 -207 -71
rect -147 -37 -89 -31
rect -147 -71 -135 -37
rect -101 -71 -89 -37
rect -147 -77 -89 -71
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect 89 -37 147 -31
rect 89 -71 101 -37
rect 135 -71 147 -37
rect 89 -77 147 -71
rect 207 -37 265 -31
rect 207 -71 219 -37
rect 253 -71 265 -37
rect 207 -77 265 -71
rect 325 -37 383 -31
rect 325 -71 337 -37
rect 371 -71 383 -37
rect 325 -77 383 -71
rect 443 -37 501 -31
rect 443 -71 455 -37
rect 489 -71 501 -37
rect 443 -77 501 -71
rect 561 -37 619 -31
rect 561 -71 573 -37
rect 607 -71 619 -37
rect 561 -77 619 -71
rect 679 -37 737 -31
rect 679 -71 691 -37
rect 725 -71 737 -37
rect 679 -77 737 -71
rect 797 -37 855 -31
rect 797 -71 809 -37
rect 843 -71 855 -37
rect 797 -77 855 -71
rect 915 -37 973 -31
rect 915 -71 927 -37
rect 961 -71 973 -37
rect 915 -77 973 -71
rect 1033 -37 1091 -31
rect 1033 -71 1045 -37
rect 1079 -71 1091 -37
rect 1033 -77 1091 -71
rect 1151 -37 1209 -31
rect 1151 -71 1163 -37
rect 1197 -71 1209 -37
rect 1151 -77 1209 -71
rect 1269 -37 1327 -31
rect 1269 -71 1281 -37
rect 1315 -71 1327 -37
rect 1269 -77 1327 -71
rect 1387 -37 1445 -31
rect 1387 -71 1399 -37
rect 1433 -71 1445 -37
rect 1387 -77 1445 -71
rect -1498 -130 -1452 -118
rect -1498 -706 -1492 -130
rect -1458 -706 -1452 -130
rect -1498 -718 -1452 -706
rect -1380 -130 -1334 -118
rect -1380 -706 -1374 -130
rect -1340 -706 -1334 -130
rect -1380 -718 -1334 -706
rect -1262 -130 -1216 -118
rect -1262 -706 -1256 -130
rect -1222 -706 -1216 -130
rect -1262 -718 -1216 -706
rect -1144 -130 -1098 -118
rect -1144 -706 -1138 -130
rect -1104 -706 -1098 -130
rect -1144 -718 -1098 -706
rect -1026 -130 -980 -118
rect -1026 -706 -1020 -130
rect -986 -706 -980 -130
rect -1026 -718 -980 -706
rect -908 -130 -862 -118
rect -908 -706 -902 -130
rect -868 -706 -862 -130
rect -908 -718 -862 -706
rect -790 -130 -744 -118
rect -790 -706 -784 -130
rect -750 -706 -744 -130
rect -790 -718 -744 -706
rect -672 -130 -626 -118
rect -672 -706 -666 -130
rect -632 -706 -626 -130
rect -672 -718 -626 -706
rect -554 -130 -508 -118
rect -554 -706 -548 -130
rect -514 -706 -508 -130
rect -554 -718 -508 -706
rect -436 -130 -390 -118
rect -436 -706 -430 -130
rect -396 -706 -390 -130
rect -436 -718 -390 -706
rect -318 -130 -272 -118
rect -318 -706 -312 -130
rect -278 -706 -272 -130
rect -318 -718 -272 -706
rect -200 -130 -154 -118
rect -200 -706 -194 -130
rect -160 -706 -154 -130
rect -200 -718 -154 -706
rect -82 -130 -36 -118
rect -82 -706 -76 -130
rect -42 -706 -36 -130
rect -82 -718 -36 -706
rect 36 -130 82 -118
rect 36 -706 42 -130
rect 76 -706 82 -130
rect 36 -718 82 -706
rect 154 -130 200 -118
rect 154 -706 160 -130
rect 194 -706 200 -130
rect 154 -718 200 -706
rect 272 -130 318 -118
rect 272 -706 278 -130
rect 312 -706 318 -130
rect 272 -718 318 -706
rect 390 -130 436 -118
rect 390 -706 396 -130
rect 430 -706 436 -130
rect 390 -718 436 -706
rect 508 -130 554 -118
rect 508 -706 514 -130
rect 548 -706 554 -130
rect 508 -718 554 -706
rect 626 -130 672 -118
rect 626 -706 632 -130
rect 666 -706 672 -130
rect 626 -718 672 -706
rect 744 -130 790 -118
rect 744 -706 750 -130
rect 784 -706 790 -130
rect 744 -718 790 -706
rect 862 -130 908 -118
rect 862 -706 868 -130
rect 902 -706 908 -130
rect 862 -718 908 -706
rect 980 -130 1026 -118
rect 980 -706 986 -130
rect 1020 -706 1026 -130
rect 980 -718 1026 -706
rect 1098 -130 1144 -118
rect 1098 -706 1104 -130
rect 1138 -706 1144 -130
rect 1098 -718 1144 -706
rect 1216 -130 1262 -118
rect 1216 -706 1222 -130
rect 1256 -706 1262 -130
rect 1216 -718 1262 -706
rect 1334 -130 1380 -118
rect 1334 -706 1340 -130
rect 1374 -706 1380 -130
rect 1334 -718 1380 -706
rect 1452 -130 1498 -118
rect 1452 -706 1458 -130
rect 1492 -706 1498 -130
rect 1452 -718 1498 -706
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -1589 -884 1589 884
string parameters w 3 l 0.3 m 2 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
