magic
tech sky130A
magscale 1 2
timestamp 1663665886
<< nwell >>
rect 7230 534660 7480 536800
rect 7230 534610 7540 534660
rect 575550 365240 575860 365290
rect 575610 363100 575860 365240
rect 578350 365240 578660 365290
rect 578410 363100 578660 365240
<< pwell >>
rect 514250 667660 514780 668110
rect 514250 665410 514790 667660
rect 514250 664950 514780 665410
rect 506460 572000 506990 572450
rect 506460 569750 507000 572000
rect 506460 569290 506990 569750
rect 559050 569420 559580 572580
rect 7900 534610 8410 536800
rect 566000 485110 569160 485640
rect 574680 363100 575190 365290
rect 577480 363100 577990 365290
rect 2970 324053 6130 324583
<< nmos >>
rect 514420 666100 514620 666500
rect 506630 570440 506830 570840
rect 559220 569980 559420 571980
rect 566560 485270 568560 485470
rect 3530 324213 5530 324413
<< ndiff >>
rect 514420 666660 514620 666700
rect 514420 666540 514460 666660
rect 514580 666540 514620 666660
rect 514420 666500 514620 666540
rect 514420 666060 514620 666100
rect 514420 665930 514450 666060
rect 514580 665930 514620 666060
rect 514420 665900 514620 665930
rect 559220 572140 559420 572180
rect 559220 572020 559260 572140
rect 559380 572020 559420 572140
rect 559220 571980 559420 572020
rect 506630 571000 506830 571040
rect 506630 570880 506670 571000
rect 506790 570880 506830 571000
rect 506630 570840 506830 570880
rect 506630 570400 506830 570440
rect 506630 570270 506660 570400
rect 506790 570270 506830 570400
rect 506630 570240 506830 570270
rect 559220 569940 559420 569980
rect 559220 569820 559260 569940
rect 559380 569820 559420 569940
rect 559220 569780 559420 569820
rect 566360 485430 566560 485470
rect 566360 485310 566400 485430
rect 566520 485310 566560 485430
rect 566360 485270 566560 485310
rect 568560 485430 568760 485470
rect 568560 485310 568600 485430
rect 568720 485310 568760 485430
rect 568560 485270 568760 485310
rect 3330 324373 3530 324413
rect 3330 324253 3370 324373
rect 3490 324253 3530 324373
rect 3330 324213 3530 324253
rect 5530 324373 5730 324413
rect 5530 324253 5570 324373
rect 5690 324253 5730 324373
rect 5530 324213 5730 324253
<< ndiffc >>
rect 514460 666540 514580 666660
rect 514450 665930 514580 666060
rect 559260 572020 559380 572140
rect 506670 570880 506790 571000
rect 506660 570270 506790 570400
rect 559260 569820 559380 569940
rect 566400 485310 566520 485430
rect 568600 485310 568720 485430
rect 3370 324253 3490 324373
rect 5570 324253 5690 324373
<< psubdiff >>
rect 514420 666860 514620 666900
rect 514420 666740 514460 666860
rect 514580 666740 514620 666860
rect 514420 666700 514620 666740
rect 559220 572340 559420 572380
rect 559220 572220 559260 572340
rect 559380 572220 559420 572340
rect 559220 572180 559420 572220
rect 506630 571200 506830 571240
rect 506630 571080 506670 571200
rect 506790 571080 506830 571200
rect 506630 571040 506830 571080
rect 8250 536730 8360 536760
rect 8250 534700 8280 536730
rect 8330 534700 8360 536730
rect 8250 534660 8360 534700
rect 568760 485430 568960 485470
rect 568760 485310 568800 485430
rect 568920 485310 568960 485430
rect 568760 485270 568960 485310
rect 574730 365200 574840 365240
rect 574730 363170 574760 365200
rect 574810 363170 574840 365200
rect 574730 363140 574840 363170
rect 577530 365200 577640 365240
rect 577530 363170 577560 365200
rect 577610 363170 577640 365200
rect 577530 363140 577640 363170
rect 5730 324373 5930 324413
rect 5730 324253 5770 324373
rect 5890 324253 5930 324373
rect 5730 324213 5930 324253
<< nsubdiff >>
rect 7270 536720 7400 536760
rect 7270 534680 7300 536720
rect 7370 534680 7400 536720
rect 7270 534660 7400 534680
rect 575690 365220 575820 365240
rect 575690 363180 575720 365220
rect 575790 363180 575820 365220
rect 575690 363140 575820 363180
rect 578490 365220 578620 365240
rect 578490 363180 578520 365220
rect 578590 363180 578620 365220
rect 578490 363140 578620 363180
<< psubdiffcont >>
rect 514460 666740 514580 666860
rect 559260 572220 559380 572340
rect 506670 571080 506790 571200
rect 8280 534700 8330 536730
rect 568800 485310 568920 485430
rect 574760 363170 574810 365200
rect 577560 363170 577610 365200
rect 5770 324253 5890 324373
<< nsubdiffcont >>
rect 7300 534680 7370 536720
rect 575720 363180 575790 365220
rect 578520 363180 578590 365220
<< poly >>
rect 514330 666100 514420 666500
rect 514620 666450 515490 666500
rect 514620 666140 515050 666450
rect 515450 666140 515490 666450
rect 514620 666100 515490 666140
rect 506540 570440 506630 570840
rect 506830 570790 507700 570840
rect 506830 570480 507260 570790
rect 507660 570480 507700 570790
rect 506830 570440 507700 570480
rect 559130 569980 559220 571980
rect 559420 571930 559810 571980
rect 559420 570030 559520 571930
rect 559760 570030 559810 571930
rect 559420 569980 559810 570030
rect 566560 485470 568560 485560
rect 566560 485170 568560 485270
rect 566560 484930 566610 485170
rect 568510 484930 568560 485170
rect 566560 484880 568560 484930
rect 3530 324413 5530 324503
rect 3530 324113 5530 324213
rect 3530 323873 3580 324113
rect 5480 323873 5530 324113
rect 3530 323823 5530 323873
<< polycont >>
rect 515050 666140 515450 666450
rect 507260 570480 507660 570790
rect 559520 570030 559760 571930
rect 566610 484930 568510 485170
rect 3580 323873 5480 324113
<< locali >>
rect 514440 667870 514600 667890
rect 514440 667570 514450 667870
rect 514440 666540 514460 667570
rect 514580 666540 514600 667870
rect 514440 666520 514600 666540
rect 514930 666450 515490 666500
rect 514930 666140 515050 666450
rect 515450 666140 515490 666450
rect 514930 666100 515490 666140
rect 514430 666060 514600 666080
rect 514430 665990 514450 666060
rect 514440 665930 514450 665990
rect 514580 665930 514600 666060
rect 514440 665890 514600 665930
rect 514440 665330 514460 665890
rect 514420 665300 514460 665330
rect 514580 665330 514600 665890
rect 514580 665300 514620 665330
rect 506650 572210 506810 572230
rect 506650 571910 506660 572210
rect 506650 570880 506670 571910
rect 506790 570880 506810 572210
rect 506650 570860 506810 570880
rect 507140 570790 507700 570840
rect 507140 570480 507260 570790
rect 507660 570480 507700 570790
rect 507140 570440 507700 570480
rect 506640 570400 506810 570420
rect 506640 570330 506660 570400
rect 506650 570270 506660 570330
rect 506790 570270 506810 570400
rect 506650 570230 506810 570270
rect 506650 569670 506670 570230
rect 506630 569640 506670 569670
rect 506790 569670 506810 570230
rect 506790 569640 506830 569670
rect 559240 572340 559400 572360
rect 559240 572040 559250 572340
rect 559240 572020 559260 572040
rect 559380 572020 559400 572340
rect 559240 572000 559400 572020
rect 559490 571930 559790 571960
rect 559490 570030 559520 571930
rect 559760 570030 559790 571930
rect 559490 570000 559790 570030
rect 559240 569940 559400 569960
rect 559240 569800 559260 569940
rect 559220 569770 559260 569800
rect 559380 569800 559400 569940
rect 559380 569770 559420 569800
rect 582200 540310 585180 555620
rect 7270 536720 7400 536760
rect 7270 534680 7300 536720
rect 7370 534680 7400 536720
rect 8260 536730 8350 536750
rect 7270 534660 7400 534680
rect 8260 534700 8280 536730
rect 8330 534700 8350 536730
rect 8260 534670 8350 534700
rect 566350 485450 566380 485470
rect 566350 485430 566540 485450
rect 566520 485310 566540 485430
rect 566350 485290 566540 485310
rect 568580 485440 568940 485450
rect 568580 485430 568620 485440
rect 568580 485310 568600 485430
rect 568920 485310 568940 485440
rect 568580 485290 568940 485310
rect 566350 485270 566380 485290
rect 566580 485170 568540 485200
rect 566580 484930 566610 485170
rect 568510 484930 568540 485170
rect 566580 484900 568540 484930
rect 574740 365200 574830 365230
rect 574740 363170 574760 365200
rect 574810 363170 574830 365200
rect 575690 365220 575820 365240
rect 574740 363150 574830 363170
rect 575690 363180 575720 365220
rect 575790 363180 575820 365220
rect 575690 363140 575820 363180
rect 577540 365200 577630 365230
rect 577540 363170 577560 365200
rect 577610 363170 577630 365200
rect 578490 365220 578620 365240
rect 577540 363150 577630 363170
rect 578490 363180 578520 365220
rect 578590 363180 578620 365220
rect 578490 363140 578620 363180
rect 3320 324393 3350 324413
rect 3320 324373 3510 324393
rect 3490 324253 3510 324373
rect 3320 324233 3510 324253
rect 5550 324383 5910 324393
rect 5550 324373 5590 324383
rect 5550 324253 5570 324373
rect 5890 324253 5910 324383
rect 5550 324233 5910 324253
rect 3320 324213 3350 324233
rect 3550 324113 5510 324143
rect 3550 323873 3580 324113
rect 5480 323873 5510 324113
rect 3550 323843 5510 323873
<< viali >>
rect 15690 701230 21540 703180
rect 67850 701700 73380 703110
rect 228670 701850 232530 702520
rect 330480 701740 334340 702410
rect 463720 699400 471140 701590
rect 510880 696600 525130 703440
rect 566440 699450 573030 701120
rect 1340 679860 3090 685550
rect 580470 678030 581910 682990
rect 498670 667090 500420 668100
rect 514450 667570 514580 667870
rect 514460 666860 514580 667570
rect 514460 666740 514580 666860
rect 514460 666660 514580 666740
rect 514460 666540 514580 666660
rect 515050 666140 515450 666450
rect 514460 665300 514580 665890
rect 514320 664830 514680 665300
rect 520580 664340 526480 669740
rect 520780 641340 526680 646740
rect 576690 630020 583530 644270
rect 520580 617740 526580 623040
rect 577730 580390 583180 583570
rect 490680 571430 492430 572440
rect 506660 571910 506790 572210
rect 506670 571200 506790 571910
rect 506670 571080 506790 571200
rect 506670 571000 506790 571080
rect 506670 570880 506790 571000
rect 507260 570480 507660 570790
rect 506670 569640 506790 570230
rect 506530 569170 506890 569640
rect 512590 568680 518490 574080
rect 543270 571560 545020 572570
rect 559250 572220 559260 572340
rect 559260 572220 559380 572340
rect 559250 572140 559380 572220
rect 559250 572040 559260 572140
rect 559260 572040 559380 572140
rect 559520 570110 559760 571840
rect 559260 569820 559380 569940
rect 559260 569770 559380 569820
rect 559120 569300 559480 569770
rect 565180 568810 571080 574210
rect 870 549250 2600 564320
rect 512790 545680 518690 551080
rect 565380 545810 571280 551210
rect 6920 534720 7200 536700
rect 7300 534680 7370 536720
rect 7830 536320 7870 536740
rect 8280 534700 8330 536730
rect 8420 534720 8700 536700
rect 512590 522080 518590 527380
rect 565180 522210 571180 527510
rect 300 511100 2350 512460
rect 568140 499670 569150 501420
rect 580590 493390 582340 495690
rect 565880 485430 566350 485570
rect 565880 485310 566400 485430
rect 566400 485310 566520 485430
rect 565880 485210 566350 485310
rect 568620 485430 568920 485440
rect 568620 485310 568720 485430
rect 568720 485310 568800 485430
rect 568800 485310 568920 485430
rect 566690 484930 568420 485170
rect 518790 473510 524090 479510
rect 542390 473410 547790 479310
rect 565390 473610 570790 479510
rect 330 467850 2380 469210
rect 576750 448670 578500 450970
rect 400 423400 1800 424600
rect 571720 405820 577750 407140
rect 400 380100 1800 381300
rect 574760 363170 574810 365200
rect 575220 363160 575260 363580
rect 575720 363180 575790 365220
rect 577560 363170 577610 365200
rect 578020 363160 578060 363580
rect 578520 363180 578590 365220
rect 579150 359440 582190 360800
rect 400 336900 1800 338100
rect 9373 329630 11123 329860
rect 9360 328850 11123 329630
rect 2850 324373 3320 324513
rect 2850 324253 3370 324373
rect 3370 324253 3490 324373
rect 2850 324153 3320 324253
rect 5590 324373 5890 324383
rect 5590 324253 5690 324373
rect 5690 324253 5770 324373
rect 5770 324253 5890 324373
rect 3660 323873 5390 324113
rect 9360 324110 11100 328850
rect 3800 322000 7400 323000
rect 400 294900 1800 296100
rect 573690 269790 579290 270990
rect 400 251800 1800 253000
rect 579460 198160 580960 201000
rect 579500 189900 580900 198160
rect 700 163110 2330 177370
rect 576400 167200 579400 175500
rect 573200 151830 576200 152000
rect 573150 148990 576200 151830
rect 573200 143700 576200 148990
rect 400 124300 1800 125500
rect 570850 123400 577320 130770
<< metal1 >>
rect 10900 703180 21970 703660
rect 10900 701470 15690 703180
rect 10890 701230 15690 701470
rect 21540 701230 21970 703180
rect 10890 700970 21970 701230
rect 930 685550 9060 685890
rect 930 679860 1340 685550
rect 3090 685420 9060 685550
rect 3090 679860 9140 685420
rect 930 679650 9140 679860
rect 330 564320 3200 564730
rect 330 549250 870 564320
rect 2600 549250 3200 564320
rect 330 548720 3200 549250
rect 8110 539100 9140 679650
rect 5640 538420 9140 539100
rect 5640 534580 6320 538420
rect 7660 536860 9860 537540
rect 7270 536740 7500 536760
rect 6880 536720 7500 536740
rect 7720 536740 7960 536860
rect 7720 536730 7830 536740
rect 6880 536700 7300 536720
rect 6880 534720 6920 536700
rect 7200 534720 7300 536700
rect 6880 534680 7300 534720
rect 7370 534680 7500 536720
rect 7800 536320 7830 536730
rect 7870 536730 7960 536740
rect 8120 536740 8350 536750
rect 8120 536730 8740 536740
rect 7870 536320 7890 536730
rect 7800 536290 7890 536320
rect 7270 534660 7500 534680
rect 7710 534790 7760 536130
rect 7710 534580 7770 534790
rect 8120 534700 8280 536730
rect 8330 536700 8740 536730
rect 8330 534720 8420 536700
rect 8700 534720 8740 536700
rect 8330 534700 8740 534720
rect 8120 534680 8740 534700
rect 8120 534670 8350 534680
rect 5640 533900 7840 534580
rect 9260 533800 9860 536860
rect 8340 533400 9900 533800
rect 8350 532720 9060 533400
rect 7170 532450 7350 532620
rect 8350 532610 8700 532720
rect 7230 531980 7370 532150
rect 7200 531950 7370 531980
rect 9610 532060 9750 532070
rect 9610 531950 9810 532060
rect 7200 531860 7340 531950
rect 9670 531940 9810 531950
rect 9630 531500 9770 531510
rect 7230 531370 7370 531490
rect 9630 531480 9800 531500
rect 9630 531390 9810 531480
rect 9660 531380 9810 531390
rect 9670 531360 9810 531380
rect 7220 530810 7360 530930
rect 9650 530110 9790 530230
rect 8120 525610 8310 527830
rect 7770 525470 8310 525610
rect 6280 525390 8310 525470
rect 6270 525270 8310 525390
rect 8510 525470 8610 527760
rect 8770 526200 8850 527650
rect 8880 526810 8960 527650
rect 10890 526810 11920 700970
rect 15390 700950 21970 700970
rect 67550 703110 73630 703460
rect 67550 701700 67850 703110
rect 73380 701700 73630 703110
rect 12950 698940 24950 698960
rect 67550 698940 73630 701700
rect 228240 702520 233100 703020
rect 228240 701850 228670 702520
rect 232530 701850 233100 702520
rect 228240 701380 233100 701850
rect 228230 701360 233100 701380
rect 330040 702850 456370 702910
rect 330040 702410 457240 702850
rect 330040 701740 330480 702410
rect 334340 701740 457240 702410
rect 228230 698980 233080 701360
rect 330040 701240 457240 701740
rect 12950 697690 73820 698940
rect 8880 526430 11920 526810
rect 8880 526390 11910 526430
rect 8880 526380 10910 526390
rect 12970 526200 14000 697690
rect 228230 696670 452570 698980
rect 455570 697640 457240 701240
rect 463060 701650 471790 703560
rect 510600 703440 525450 703780
rect 463060 701590 506390 701650
rect 463060 699400 463720 701590
rect 471140 699400 506390 701590
rect 463060 698690 506390 699400
rect 469180 698670 506390 698690
rect 498560 697640 500610 697700
rect 228330 696640 452570 696670
rect 450030 694770 452570 696640
rect 455440 695970 500620 697640
rect 450030 694750 497150 694770
rect 450030 693100 497500 694750
rect 450030 692770 452570 693100
rect 495510 674560 497500 693100
rect 498560 692400 500610 695970
rect 503600 694930 506390 698670
rect 510600 696600 510880 703440
rect 525130 696600 525450 703440
rect 510600 696230 525450 696600
rect 566000 701120 573590 702930
rect 566000 699450 566440 701120
rect 573030 699450 573590 701120
rect 566000 695050 573590 699450
rect 503600 693460 563610 694930
rect 503600 692670 563660 693460
rect 503600 692640 506390 692670
rect 495540 666500 497500 674560
rect 498570 674210 500560 692400
rect 561240 684580 563660 692670
rect 498570 668100 500530 674210
rect 498570 667090 498670 668100
rect 500420 667090 500530 668100
rect 519680 669740 527080 670340
rect 495640 665560 497460 666500
rect 498570 666470 500530 667090
rect 514270 667870 514760 668060
rect 514270 667570 514450 667870
rect 514580 667650 514760 667870
rect 495640 665530 497440 665560
rect 497280 664200 497420 665530
rect 498600 665490 500530 666470
rect 501760 666940 503720 666960
rect 501760 666140 506880 666940
rect 514270 666540 514460 667570
rect 514580 666540 514790 667650
rect 519680 667400 520580 669740
rect 514270 666530 514790 666540
rect 514420 666500 514620 666530
rect 515020 666450 520580 667400
rect 515020 666140 515050 666450
rect 515450 666140 520580 666450
rect 501760 665770 506980 666140
rect 514420 666070 514620 666100
rect 501780 665640 506980 665770
rect 501780 665580 503710 665640
rect 498640 665480 500510 665490
rect 498640 664280 498780 665480
rect 497620 663960 498780 664280
rect 501780 664210 502230 665580
rect 505480 658440 506980 665640
rect 514270 665890 514760 666070
rect 514270 665300 514460 665890
rect 514580 665300 514760 665890
rect 515020 665600 520580 666140
rect 514270 664960 514320 665300
rect 514280 664830 514320 664960
rect 514680 664830 514760 665300
rect 514280 664800 514760 664830
rect 519680 664340 520580 665600
rect 526480 664340 527080 669740
rect 519680 663640 527080 664340
rect 505480 657140 514480 658440
rect 503450 653460 503690 653490
rect 503450 652270 503480 653460
rect 503670 652270 503690 653460
rect 503450 652240 503690 652270
rect 512880 645040 514380 657140
rect 519780 646740 527180 647440
rect 519780 645040 520780 646740
rect 512880 642440 520780 645040
rect 514380 642340 520780 642440
rect 519780 641340 520780 642340
rect 526680 641340 527180 646740
rect 519780 640740 527180 641340
rect 519880 623040 527180 623740
rect 519880 617740 520580 623040
rect 526580 617740 527180 623040
rect 519880 617040 527180 617740
rect 487540 598170 493100 598200
rect 561300 598170 563600 684580
rect 487540 596830 563600 598170
rect 487520 595370 563600 596830
rect 487520 595230 563590 595370
rect 487520 595190 493100 595230
rect 487520 582420 489540 595190
rect 567180 592420 569480 695050
rect 571390 683050 583580 683560
rect 571370 682990 583580 683050
rect 571370 680010 580470 682990
rect 571390 678030 580470 680010
rect 581910 678030 583580 682990
rect 571390 677700 583580 678030
rect 491720 592400 569520 592420
rect 490590 589480 569520 592400
rect 487550 570840 489510 582420
rect 490590 582130 493070 589480
rect 567180 589370 569480 589480
rect 571400 587910 573510 677700
rect 576350 644270 583900 644590
rect 576350 630020 576690 644270
rect 583530 630020 583900 644270
rect 576350 629740 583900 630020
rect 547990 587880 573510 587910
rect 540120 584500 573510 587880
rect 490590 582110 493120 582130
rect 490580 579750 493120 582110
rect 490580 572440 492540 579750
rect 490580 571430 490680 572440
rect 492430 571430 492540 572440
rect 511690 574080 519090 574680
rect 487650 569900 489470 570840
rect 490580 570810 492540 571430
rect 506480 572210 506970 572400
rect 506480 571910 506660 572210
rect 506790 571990 506970 572210
rect 487650 569870 489450 569900
rect 489290 568540 489430 569870
rect 490610 569830 492540 570810
rect 493770 571280 495730 571300
rect 493770 570480 498890 571280
rect 506480 570880 506670 571910
rect 506790 570880 507000 571990
rect 511690 571740 512590 574080
rect 506480 570870 507000 570880
rect 506630 570840 506830 570870
rect 507230 570790 512590 571740
rect 507230 570480 507260 570790
rect 507660 570480 512590 570790
rect 493770 570110 498990 570480
rect 506630 570410 506830 570440
rect 493790 569980 498990 570110
rect 493790 569920 495720 569980
rect 490650 569820 492520 569830
rect 490650 568620 490790 569820
rect 489630 568300 490790 568620
rect 493790 568550 494240 569920
rect 497490 562780 498990 569980
rect 506480 570230 506970 570410
rect 506480 569640 506670 570230
rect 506790 569640 506970 570230
rect 507230 569940 512590 570480
rect 506480 569300 506530 569640
rect 506490 569170 506530 569300
rect 506890 569170 506970 569640
rect 506490 569140 506970 569170
rect 511690 568680 512590 569940
rect 518490 568680 519090 574080
rect 540140 570970 542100 584500
rect 547990 584480 573510 584500
rect 577270 583570 583810 584240
rect 577270 582260 577730 583570
rect 543280 582240 577730 582260
rect 543170 580390 577730 582240
rect 583180 580390 583810 583570
rect 543170 579880 583810 580390
rect 543170 572570 545130 579880
rect 577270 579860 583810 579880
rect 543170 571560 543270 572570
rect 545020 571560 545130 572570
rect 564280 574210 571680 574810
rect 559070 572340 559560 572530
rect 559070 572040 559250 572340
rect 559380 572040 559560 572340
rect 559070 572000 559560 572040
rect 564280 571870 565180 574210
rect 540240 570030 542060 570970
rect 543170 570940 545130 571560
rect 559490 571840 565180 571870
rect 540240 570000 542040 570030
rect 511690 567980 519090 568680
rect 541880 568670 542020 570000
rect 543200 569960 545130 570940
rect 546360 571410 548320 571430
rect 546360 570610 551480 571410
rect 546360 570240 551580 570610
rect 546380 570110 551580 570240
rect 546380 570050 548310 570110
rect 543240 569950 545110 569960
rect 543240 568750 543380 569950
rect 542220 568430 543380 568750
rect 546380 568680 546830 570050
rect 550080 562910 551580 570110
rect 559490 570110 559520 571840
rect 559760 570110 565180 571840
rect 559490 570070 565180 570110
rect 559070 569940 559560 569960
rect 559070 569770 559260 569940
rect 559380 569770 559560 569940
rect 559070 569430 559120 569770
rect 559080 569300 559120 569430
rect 559480 569300 559560 569770
rect 559080 569270 559560 569300
rect 564280 568810 565180 570070
rect 571080 568810 571680 574210
rect 564280 568110 571680 568810
rect 497490 561480 506490 562780
rect 550080 561610 559080 562910
rect 495460 557800 495700 557830
rect 495460 556610 495490 557800
rect 495680 556610 495700 557800
rect 495460 556580 495700 556610
rect 504890 549380 506390 561480
rect 548050 557930 548290 557960
rect 548050 556740 548080 557930
rect 548270 556740 548290 557930
rect 548050 556710 548290 556740
rect 511790 551080 519190 551780
rect 511790 549380 512790 551080
rect 504890 546780 512790 549380
rect 506390 546680 512790 546780
rect 511790 545680 512790 546680
rect 518690 545680 519190 551080
rect 557480 549510 558980 561610
rect 564380 551210 571780 551910
rect 564380 549510 565380 551210
rect 557480 546910 565380 549510
rect 558980 546810 565380 546910
rect 511790 545080 519190 545680
rect 564380 545810 565380 546810
rect 571280 545810 571780 551210
rect 564380 545210 571780 545810
rect 511890 527380 519190 528080
rect 8770 525780 14010 526200
rect 6270 512620 7290 525270
rect 8510 524980 9520 525470
rect 130 512460 7290 512620
rect 130 511100 300 512460
rect 2350 511100 7290 512460
rect 130 510940 7290 511100
rect 8490 524430 9520 524980
rect 130 510930 5960 510940
rect 8490 469370 9510 524430
rect 511890 522080 512590 527380
rect 518590 522080 519190 527380
rect 511890 521380 519190 522080
rect 564480 527510 571780 528210
rect 564480 522210 565180 527510
rect 571180 522210 571780 527510
rect 564480 521510 571780 522210
rect 567550 504450 582650 504550
rect 566580 504130 582650 504450
rect 566580 502810 582680 504130
rect 565250 502670 582680 502810
rect 566580 502650 582680 502670
rect 566610 502630 582680 502650
rect 567550 502590 582680 502630
rect 565010 501450 565330 502470
rect 567520 501490 578820 501520
rect 566540 501450 578820 501490
rect 565010 501420 578820 501450
rect 565010 501310 568140 501420
rect 566530 499670 568140 501310
rect 569150 501410 578820 501420
rect 569150 499670 578840 501410
rect 566530 499580 578840 499670
rect 566540 499560 578840 499580
rect 566820 498310 568010 498330
rect 565260 497860 568010 498310
rect 553290 496610 554540 496640
rect 553290 496420 553320 496610
rect 554510 496420 554540 496610
rect 553290 496400 554540 496420
rect 566630 496380 568010 497860
rect 566690 496370 568010 496380
rect 566690 494610 567990 496370
rect 558190 493210 567990 494610
rect 558190 493110 567190 493210
rect 558190 487210 559490 493110
rect 543490 485710 559490 487210
rect 543390 480310 546090 485710
rect 558190 485610 559490 485710
rect 566010 485610 566540 485620
rect 565850 485570 566540 485610
rect 565850 485210 565880 485570
rect 566350 485430 566540 485570
rect 566520 485310 566540 485430
rect 566350 485210 566540 485310
rect 565850 485130 566540 485210
rect 568580 485440 569110 485620
rect 568580 485310 568620 485440
rect 568920 485310 569110 485440
rect 566650 485170 568450 485200
rect 566650 484930 566690 485170
rect 568420 484930 568450 485170
rect 568580 485130 569110 485310
rect 566650 480410 568450 484930
rect 518090 479510 524790 480210
rect 518090 473510 518790 479510
rect 524090 473510 524790 479510
rect 518090 472910 524790 473510
rect 541790 479310 548490 480310
rect 541790 473410 542390 479310
rect 547790 473410 548490 479310
rect 541790 472910 548490 473410
rect 564690 479510 571390 480410
rect 564690 473610 565390 479510
rect 570790 473610 571390 479510
rect 564690 473010 571390 473610
rect 180 469210 9510 469370
rect 180 467850 330 469210
rect 2380 467850 9510 469210
rect 180 467700 9510 467850
rect 8490 467680 9510 467700
rect 576460 450970 578840 499560
rect 580300 495690 582680 502590
rect 580300 493390 580590 495690
rect 582340 493390 582680 495690
rect 580300 493190 582680 493390
rect 576460 448670 576750 450970
rect 578500 448670 578840 450970
rect 576460 448470 578840 448670
rect 200 424600 2000 424800
rect 200 423400 400 424600
rect 1800 423400 2000 424600
rect 200 423200 2000 423400
rect 571340 407350 575660 408050
rect 571340 407140 583800 407350
rect 571340 405820 571720 407140
rect 577750 405820 583800 407140
rect 571340 405610 583800 405820
rect 200 381300 2000 381500
rect 200 380100 400 381300
rect 1800 380100 2000 381300
rect 200 379900 2000 380100
rect 571340 366400 575660 405610
rect 578050 366600 582350 366740
rect 571340 365400 575800 366400
rect 577800 365800 582350 366600
rect 577800 365400 578200 365800
rect 571340 365300 572780 365400
rect 574740 365200 574970 365230
rect 574740 365000 574760 365200
rect 573800 364800 574760 365000
rect 573800 363400 574000 364800
rect 574600 363400 574760 364800
rect 573800 363200 574760 363400
rect 574740 363170 574760 363200
rect 574810 363170 574970 365200
rect 575320 365110 575380 365400
rect 575330 363770 575380 365110
rect 575590 365220 575820 365240
rect 574740 363150 574970 363170
rect 575200 363580 575290 363610
rect 575200 363160 575220 363580
rect 575260 363160 575290 363580
rect 575200 362880 575290 363160
rect 575590 363180 575720 365220
rect 575790 365200 575820 365220
rect 577540 365200 577770 365230
rect 575790 365000 576200 365200
rect 577540 365000 577560 365200
rect 575790 363400 575800 365000
rect 576000 363400 576200 365000
rect 575790 363200 576200 363400
rect 576600 364800 577560 365000
rect 576600 363400 576800 364800
rect 577400 363400 577560 364800
rect 576600 363200 577560 363400
rect 575790 363180 575820 363200
rect 575590 363140 575820 363180
rect 577540 363170 577560 363200
rect 577610 363170 577770 365200
rect 578120 365190 578220 365400
rect 578390 365220 578620 365240
rect 578120 365110 578180 365190
rect 578130 363770 578180 365110
rect 577540 363150 577770 363170
rect 578000 363580 578090 363610
rect 578000 363160 578020 363580
rect 578060 363160 578090 363580
rect 578000 363120 578090 363160
rect 578390 363180 578520 365220
rect 578590 365200 578620 365220
rect 578590 365000 579000 365200
rect 578590 363400 578600 365000
rect 578800 363400 579000 365000
rect 578590 363200 579000 363400
rect 578590 363180 578620 363200
rect 578390 363140 578620 363180
rect 577990 362960 578090 363120
rect 577990 362880 578110 362960
rect 575200 362240 576570 362880
rect 575630 361610 576570 362240
rect 576670 362240 578110 362880
rect 579400 362400 582350 365800
rect 576670 361510 577730 362240
rect 577530 361480 577730 361510
rect 579010 360900 582350 362400
rect 579010 360800 583790 360900
rect 579010 359440 579150 360800
rect 582190 359440 583790 360800
rect 579010 359300 583790 359440
rect 579010 357690 582350 359300
rect 576030 354520 576200 354540
rect 576030 354460 576050 354520
rect 576180 354460 576200 354520
rect 576030 354440 576200 354460
rect 577160 354530 577330 354550
rect 577160 354450 577180 354530
rect 577310 354450 577330 354530
rect 577160 354440 577330 354450
rect 6103 344680 6343 344710
rect 6103 343490 6123 344680
rect 6313 343490 6343 344680
rect 6103 343460 6343 343490
rect 200 338100 4313 338300
rect 200 336900 400 338100
rect 1800 336900 4313 338100
rect 200 336700 4313 336900
rect 2813 331310 4313 336700
rect 7563 331370 8013 332740
rect 11013 332670 12173 332990
rect 11013 331470 11153 332670
rect 9283 331460 11153 331470
rect 6083 331310 8013 331370
rect 2813 331180 8013 331310
rect 2813 330810 8033 331180
rect 2913 330010 8033 330810
rect 6073 329990 8033 330010
rect 9263 330480 11193 331460
rect 12373 331420 12513 332750
rect 12353 331390 14153 331420
rect 9263 330040 11223 330480
rect 12333 330450 14153 331390
rect 9263 329860 11240 330040
rect 9263 329630 9373 329860
rect 2980 324553 3510 324563
rect 2820 324513 3510 324553
rect 2820 324153 2850 324513
rect 3320 324373 3510 324513
rect 3490 324253 3510 324373
rect 3320 324153 3510 324253
rect 2820 324073 3510 324153
rect 5550 324383 6080 324563
rect 5550 324253 5590 324383
rect 5890 324253 6080 324383
rect 3620 324113 5420 324143
rect 3620 323873 3660 324113
rect 5390 323873 5420 324113
rect 5550 324073 6080 324253
rect 9263 324110 9360 329630
rect 11123 328850 11240 329860
rect 11100 324110 11240 328850
rect 3620 323200 5420 323873
rect 9263 323850 11240 324110
rect 3600 323000 7600 323200
rect 3600 322000 3800 323000
rect 7400 322000 7600 323000
rect 9263 322700 11223 323850
rect 3600 321800 7600 322000
rect 8900 296300 11300 322700
rect 12293 322000 14253 330450
rect 200 296100 11300 296300
rect 200 294900 400 296100
rect 1800 294900 11300 296100
rect 200 294700 11300 294900
rect 12200 253200 14600 322000
rect 576860 315490 579860 316870
rect 576860 314100 576980 315490
rect 579620 314100 579860 315490
rect 576860 312370 579860 314100
rect 573510 270990 583830 271200
rect 573510 269790 573690 270990
rect 579290 269790 583830 270990
rect 573510 269620 583830 269790
rect 200 253000 14600 253200
rect 200 251800 400 253000
rect 1800 251800 14600 253000
rect 200 251600 14600 251800
rect 572020 217610 572260 217640
rect 572020 216420 572040 217610
rect 572230 216420 572260 217610
rect 572020 216390 572260 216420
rect 574530 204300 574980 205670
rect 577980 205600 579140 205920
rect 577980 204400 578120 205600
rect 576250 204390 578120 204400
rect 573050 204110 574980 204300
rect 573040 181390 575000 204110
rect 576230 202480 578160 204390
rect 579340 204350 579480 205680
rect 579320 204320 581120 204350
rect 579300 204300 581120 204320
rect 400 177370 2740 177720
rect 400 163110 700 177370
rect 2330 163110 2740 177370
rect 573040 177280 575020 181390
rect 400 162870 2740 163110
rect 573060 152630 575020 177280
rect 576230 175800 578150 202480
rect 579300 201200 581200 204300
rect 579200 201000 581200 201200
rect 579200 198160 579460 201000
rect 580960 198160 581200 201000
rect 579200 189900 579500 198160
rect 580900 189900 581200 198160
rect 579200 189500 581200 189900
rect 576200 175500 579600 175800
rect 576200 167200 576400 175500
rect 579400 167200 579600 175500
rect 576200 166600 579600 167200
rect 572960 152600 575020 152630
rect 572900 152000 576700 152600
rect 572900 151830 573200 152000
rect 572900 148990 573150 151830
rect 572900 143700 573200 148990
rect 576200 143700 576700 152000
rect 572900 143300 576700 143700
rect 570290 130770 578040 131480
rect 200 125500 2000 125700
rect 200 124300 400 125500
rect 1800 124300 2000 125500
rect 200 124100 2000 124300
rect 570290 123400 570850 130770
rect 577320 123400 578040 130770
rect 570290 123020 578040 123400
<< via1 >>
rect 15690 701230 21540 703180
rect 1340 679860 3090 685550
rect 6920 534720 7200 536700
rect 8420 534720 8700 536700
rect 67850 701700 73380 703110
rect 228670 701850 232530 702520
rect 330480 701740 334340 702410
rect 463720 699400 471140 701590
rect 510880 696600 525130 703440
rect 566440 699450 573030 701120
rect 498670 667090 500420 668100
rect 514320 664830 514680 665300
rect 520580 664340 526480 669740
rect 503480 652270 503670 653460
rect 520780 641340 526680 646740
rect 520580 617740 526580 623040
rect 580470 678030 581910 682990
rect 576690 630020 583530 644270
rect 490680 571430 492430 572440
rect 506530 569170 506890 569640
rect 512590 568680 518490 574080
rect 577730 580390 583180 583570
rect 543270 571560 545020 572570
rect 559120 569300 559480 569770
rect 565180 568810 571080 574210
rect 495490 556610 495680 557800
rect 548080 556740 548270 557930
rect 512790 545680 518690 551080
rect 565380 545810 571280 551210
rect 300 511100 2350 512460
rect 512590 522080 518590 527380
rect 565180 522210 571180 527510
rect 568140 499670 569150 501420
rect 553320 496420 554510 496610
rect 565880 485210 566350 485570
rect 518790 473510 524090 479510
rect 542390 473410 547790 479310
rect 565390 473610 570790 479510
rect 330 467850 2380 469210
rect 580590 493390 582340 495690
rect 576750 448670 578500 450970
rect 400 423400 1800 424600
rect 571720 405820 577750 407140
rect 400 380100 1800 381300
rect 574000 363400 574600 364800
rect 575800 363400 576000 365000
rect 576800 363400 577400 364800
rect 578600 363400 578800 365000
rect 579150 359440 582190 360800
rect 576050 354460 576180 354520
rect 577180 354450 577310 354530
rect 6123 343490 6313 344680
rect 400 336900 1800 338100
rect 9373 329630 11123 329860
rect 2850 324153 3320 324513
rect 9360 328850 11123 329630
rect 9360 324110 11100 328850
rect 3800 322000 7400 323000
rect 400 294900 1800 296100
rect 576980 314100 579620 315490
rect 573690 269790 579290 270990
rect 400 251800 1800 253000
rect 572040 216420 572230 217610
rect 700 163110 2330 177370
rect 579460 198160 580960 201000
rect 579500 189900 580900 198160
rect 576400 167200 579400 175500
rect 573200 151830 576200 152000
rect 573150 148990 576200 151830
rect 573200 143700 576200 148990
rect 400 124300 1800 125500
rect 570850 123400 577320 130770
<< metal2 >>
rect 15390 703180 21970 703660
rect 15390 701230 15690 703180
rect 21540 701230 21970 703180
rect 67560 703110 73630 703470
rect 67560 701700 67850 703110
rect 73380 701700 73630 703110
rect 67560 701540 73630 701700
rect 228240 702520 233090 702990
rect 228240 701850 228670 702520
rect 232530 701850 233090 702520
rect 228240 701380 233090 701850
rect 330050 702410 334900 702880
rect 330050 701740 330480 702410
rect 334340 701740 334900 702410
rect 330050 701270 334900 701740
rect 463110 701590 471840 703610
rect 15390 700950 21970 701230
rect 463110 699400 463720 701590
rect 471140 699400 471840 701590
rect 510600 703440 525450 703780
rect 510600 700600 510880 703440
rect 463110 698980 471840 699400
rect 510000 696600 510880 700600
rect 525130 700600 525450 703440
rect 565960 701120 573480 702930
rect 525130 696600 526600 700600
rect 565960 699450 566440 701120
rect 573030 699450 573480 701120
rect 565960 698710 573480 699450
rect 510000 693800 526600 696600
rect 4400 693000 526600 693800
rect 4400 691600 5400 693000
rect 7000 691600 9200 693000
rect 10800 691600 14000 693000
rect 15600 691600 17000 693000
rect 18600 691600 20000 693000
rect 21600 691600 23000 693000
rect 24600 691600 26000 693000
rect 27600 691600 29000 693000
rect 30600 691600 32000 693000
rect 33600 691600 35000 693000
rect 36600 691600 38000 693000
rect 39600 691600 41000 693000
rect 42600 691600 44000 693000
rect 45600 691600 47000 693000
rect 48600 691600 50000 693000
rect 51600 691600 53000 693000
rect 54600 691600 56000 693000
rect 57600 691600 59000 693000
rect 60600 691600 62000 693000
rect 63600 691600 65000 693000
rect 66600 691600 68000 693000
rect 69600 691600 71000 693000
rect 72600 691600 74000 693000
rect 75600 691600 77000 693000
rect 78600 691600 80000 693000
rect 81600 691600 83000 693000
rect 84600 691600 86000 693000
rect 87600 691600 89000 693000
rect 90600 691600 92000 693000
rect 93600 691600 95000 693000
rect 96600 691600 98000 693000
rect 99600 691600 101000 693000
rect 102600 691600 104000 693000
rect 105600 691600 107000 693000
rect 108600 691600 110000 693000
rect 111600 691600 113000 693000
rect 114600 691600 116000 693000
rect 117600 691600 119000 693000
rect 120600 691600 122000 693000
rect 123600 691600 125000 693000
rect 126600 691600 128000 693000
rect 129600 691600 131000 693000
rect 132600 691600 134000 693000
rect 135600 691600 137000 693000
rect 138600 691600 140000 693000
rect 141600 691600 143000 693000
rect 144600 691600 146000 693000
rect 147600 691600 149000 693000
rect 150600 691600 152000 693000
rect 153600 691600 155000 693000
rect 156600 691600 158000 693000
rect 159600 691600 161000 693000
rect 162600 691600 164000 693000
rect 165600 691600 167000 693000
rect 168600 691600 170000 693000
rect 171600 691600 173000 693000
rect 174600 691600 176000 693000
rect 177600 691600 179000 693000
rect 180600 691600 182000 693000
rect 183600 691600 185000 693000
rect 186600 691600 188000 693000
rect 189600 691600 191000 693000
rect 192600 691600 194000 693000
rect 195600 691600 197000 693000
rect 198600 691600 200000 693000
rect 201600 691600 203000 693000
rect 204600 691600 206000 693000
rect 207600 691600 209000 693000
rect 210600 691600 212000 693000
rect 213600 691600 215000 693000
rect 216600 691600 218000 693000
rect 219600 691600 221000 693000
rect 222600 691600 224000 693000
rect 225600 691600 227000 693000
rect 228600 691600 230000 693000
rect 231600 691600 233000 693000
rect 234600 691600 236000 693000
rect 237600 691600 239000 693000
rect 240600 691600 242000 693000
rect 243600 691600 245000 693000
rect 246600 691600 248000 693000
rect 249600 691600 251000 693000
rect 252600 691600 254000 693000
rect 255600 691600 257000 693000
rect 258600 691600 260000 693000
rect 261600 691600 263000 693000
rect 264600 691600 266000 693000
rect 267600 691600 269000 693000
rect 270600 691600 272000 693000
rect 273600 691600 275000 693000
rect 276600 691600 278000 693000
rect 279600 691600 281000 693000
rect 282600 691600 284000 693000
rect 285600 691600 287000 693000
rect 288600 691600 290000 693000
rect 291600 691600 293000 693000
rect 294600 691600 296000 693000
rect 297600 691600 299000 693000
rect 300600 691600 302000 693000
rect 303600 691600 305000 693000
rect 306600 691600 308000 693000
rect 309600 691600 311000 693000
rect 312600 691600 314000 693000
rect 315600 691600 317000 693000
rect 318600 691600 320000 693000
rect 321600 691600 323000 693000
rect 324600 691600 326000 693000
rect 327600 691600 329000 693000
rect 330600 691600 332000 693000
rect 333600 691600 335000 693000
rect 336600 691600 338000 693000
rect 339600 691600 341000 693000
rect 342600 691600 344000 693000
rect 345600 691600 347000 693000
rect 348600 691600 350000 693000
rect 351600 691600 353000 693000
rect 354600 691600 356000 693000
rect 357600 691600 359000 693000
rect 360600 691600 362000 693000
rect 363600 691600 365000 693000
rect 366600 691600 368000 693000
rect 369600 691600 371000 693000
rect 372600 691600 374000 693000
rect 375600 691600 377000 693000
rect 378600 691600 380000 693000
rect 381600 691600 383000 693000
rect 384600 691600 386000 693000
rect 387600 691600 389000 693000
rect 390600 691600 392000 693000
rect 393600 691600 395000 693000
rect 396600 691600 398000 693000
rect 399600 691600 401000 693000
rect 402600 691600 404000 693000
rect 405600 691600 407000 693000
rect 408600 691600 410000 693000
rect 411600 691600 413000 693000
rect 414600 691600 416000 693000
rect 417600 691600 419000 693000
rect 420600 691600 422000 693000
rect 423600 691600 425000 693000
rect 426600 691600 428000 693000
rect 429600 691600 431000 693000
rect 432600 691600 434000 693000
rect 435600 691600 437000 693000
rect 438600 691600 440000 693000
rect 441600 691600 443000 693000
rect 444600 691600 446000 693000
rect 447600 691600 449000 693000
rect 450600 691600 452000 693000
rect 453600 691600 455000 693000
rect 456600 691600 458000 693000
rect 459600 691600 461000 693000
rect 462600 691600 464000 693000
rect 465600 691600 467000 693000
rect 468600 691600 470000 693000
rect 471600 691600 473000 693000
rect 474600 691600 476000 693000
rect 477600 691600 479000 693000
rect 480600 691600 482000 693000
rect 483600 691600 485000 693000
rect 486600 691600 488000 693000
rect 489600 691600 491000 693000
rect 492600 691600 494000 693000
rect 495600 691600 497000 693000
rect 498600 691600 500000 693000
rect 501600 691600 503000 693000
rect 504600 691600 506000 693000
rect 507600 691600 509000 693000
rect 510600 691600 512000 693000
rect 513600 691600 515000 693000
rect 516600 691600 518000 693000
rect 519600 691600 521000 693000
rect 522600 691600 524000 693000
rect 525600 691600 526600 693000
rect 4400 690000 526600 691600
rect 4400 688600 5400 690000
rect 7000 688600 9200 690000
rect 10800 688600 14000 690000
rect 15600 688600 17000 690000
rect 18600 688600 20000 690000
rect 21600 688600 23000 690000
rect 24600 688600 26000 690000
rect 27600 688600 29000 690000
rect 30600 688600 32000 690000
rect 33600 688600 35000 690000
rect 36600 688600 38000 690000
rect 39600 688600 41000 690000
rect 42600 688600 44000 690000
rect 45600 688600 47000 690000
rect 48600 688600 50000 690000
rect 51600 688600 53000 690000
rect 54600 688600 56000 690000
rect 57600 688600 59000 690000
rect 60600 688600 62000 690000
rect 63600 688600 65000 690000
rect 66600 688600 68000 690000
rect 69600 688600 71000 690000
rect 72600 688600 74000 690000
rect 75600 688600 77000 690000
rect 78600 688600 80000 690000
rect 81600 688600 83000 690000
rect 84600 688600 86000 690000
rect 87600 688600 89000 690000
rect 90600 688600 92000 690000
rect 93600 688600 95000 690000
rect 96600 688600 98000 690000
rect 99600 688600 101000 690000
rect 102600 688600 104000 690000
rect 105600 688600 107000 690000
rect 108600 688600 110000 690000
rect 111600 688600 113000 690000
rect 114600 688600 116000 690000
rect 117600 688600 119000 690000
rect 120600 688600 122000 690000
rect 123600 688600 125000 690000
rect 126600 688600 128000 690000
rect 129600 688600 131000 690000
rect 132600 688600 134000 690000
rect 135600 688600 137000 690000
rect 138600 688600 140000 690000
rect 141600 688600 143000 690000
rect 144600 688600 146000 690000
rect 147600 688600 149000 690000
rect 150600 688600 152000 690000
rect 153600 688600 155000 690000
rect 156600 688600 158000 690000
rect 159600 688600 161000 690000
rect 162600 688600 164000 690000
rect 165600 688600 167000 690000
rect 168600 688600 170000 690000
rect 171600 688600 173000 690000
rect 174600 688600 176000 690000
rect 177600 688600 179000 690000
rect 180600 688600 182000 690000
rect 183600 688600 185000 690000
rect 186600 688600 188000 690000
rect 189600 688600 191000 690000
rect 192600 688600 194000 690000
rect 195600 688600 197000 690000
rect 198600 688600 200000 690000
rect 201600 688600 203000 690000
rect 204600 688600 206000 690000
rect 207600 688600 209000 690000
rect 210600 688600 212000 690000
rect 213600 688600 215000 690000
rect 216600 688600 218000 690000
rect 219600 688600 221000 690000
rect 222600 688600 224000 690000
rect 225600 688600 227000 690000
rect 228600 688600 230000 690000
rect 231600 688600 233000 690000
rect 234600 688600 236000 690000
rect 237600 688600 239000 690000
rect 240600 688600 242000 690000
rect 243600 688600 245000 690000
rect 246600 688600 248000 690000
rect 249600 688600 251000 690000
rect 252600 688600 254000 690000
rect 255600 688600 257000 690000
rect 258600 688600 260000 690000
rect 261600 688600 263000 690000
rect 264600 688600 266000 690000
rect 267600 688600 269000 690000
rect 270600 688600 272000 690000
rect 273600 688600 275000 690000
rect 276600 688600 278000 690000
rect 279600 688600 281000 690000
rect 282600 688600 284000 690000
rect 285600 688600 287000 690000
rect 288600 688600 290000 690000
rect 291600 688600 293000 690000
rect 294600 688600 296000 690000
rect 297600 688600 299000 690000
rect 300600 688600 302000 690000
rect 303600 688600 305000 690000
rect 306600 688600 308000 690000
rect 309600 688600 311000 690000
rect 312600 688600 314000 690000
rect 315600 688600 317000 690000
rect 318600 688600 320000 690000
rect 321600 688600 323000 690000
rect 324600 688600 326000 690000
rect 327600 688600 329000 690000
rect 330600 688600 332000 690000
rect 333600 688600 335000 690000
rect 336600 688600 338000 690000
rect 339600 688600 341000 690000
rect 342600 688600 344000 690000
rect 345600 688600 347000 690000
rect 348600 688600 350000 690000
rect 351600 688600 353000 690000
rect 354600 688600 356000 690000
rect 357600 688600 359000 690000
rect 360600 688600 362000 690000
rect 363600 688600 365000 690000
rect 366600 688600 368000 690000
rect 369600 688600 371000 690000
rect 372600 688600 374000 690000
rect 375600 688600 377000 690000
rect 378600 688600 380000 690000
rect 381600 688600 383000 690000
rect 384600 688600 386000 690000
rect 387600 688600 389000 690000
rect 390600 688600 392000 690000
rect 393600 688600 395000 690000
rect 396600 688600 398000 690000
rect 399600 688600 401000 690000
rect 402600 688600 404000 690000
rect 405600 688600 407000 690000
rect 408600 688600 410000 690000
rect 411600 688600 413000 690000
rect 414600 688600 416000 690000
rect 417600 688600 419000 690000
rect 420600 688600 422000 690000
rect 423600 688600 425000 690000
rect 426600 688600 428000 690000
rect 429600 688600 431000 690000
rect 432600 688600 434000 690000
rect 435600 688600 437000 690000
rect 438600 688600 440000 690000
rect 441600 688600 443000 690000
rect 444600 688600 446000 690000
rect 447600 688600 449000 690000
rect 450600 688600 452000 690000
rect 453600 688600 455000 690000
rect 456600 688600 458000 690000
rect 459600 688600 461000 690000
rect 462600 688600 464000 690000
rect 465600 688600 467000 690000
rect 468600 688600 470000 690000
rect 471600 688600 473000 690000
rect 474600 688600 476000 690000
rect 477600 688600 479000 690000
rect 480600 688600 482000 690000
rect 483600 688600 485000 690000
rect 486600 688600 488000 690000
rect 489600 688600 491000 690000
rect 492600 688600 494000 690000
rect 495600 688600 497000 690000
rect 498600 688600 500000 690000
rect 501600 688600 503000 690000
rect 504600 688600 506000 690000
rect 507600 688600 509000 690000
rect 510600 688600 512000 690000
rect 513600 688600 515000 690000
rect 516600 688600 518000 690000
rect 519600 688600 521000 690000
rect 522600 688600 524000 690000
rect 525600 688600 526600 690000
rect 4400 687000 526600 688600
rect 930 685550 3360 685890
rect 930 679860 1340 685550
rect 3090 679860 3360 685550
rect 930 679660 3360 679860
rect 4400 685600 5400 687000
rect 7000 685600 9200 687000
rect 10800 685600 14000 687000
rect 15600 685600 17000 687000
rect 18600 685600 20000 687000
rect 21600 685600 23000 687000
rect 24600 685600 26000 687000
rect 27600 685600 29000 687000
rect 30600 685600 32000 687000
rect 33600 685600 35000 687000
rect 36600 685600 38000 687000
rect 39600 685600 41000 687000
rect 42600 685600 44000 687000
rect 45600 685600 47000 687000
rect 48600 685600 50000 687000
rect 51600 685600 53000 687000
rect 54600 685600 56000 687000
rect 57600 685600 59000 687000
rect 60600 685600 62000 687000
rect 63600 685600 65000 687000
rect 66600 685600 68000 687000
rect 69600 685600 71000 687000
rect 72600 685600 74000 687000
rect 75600 685600 77000 687000
rect 78600 685600 80000 687000
rect 81600 685600 83000 687000
rect 84600 685600 86000 687000
rect 87600 685600 89000 687000
rect 90600 685600 92000 687000
rect 93600 685600 95000 687000
rect 96600 685600 98000 687000
rect 99600 685600 101000 687000
rect 102600 685600 104000 687000
rect 105600 685600 107000 687000
rect 108600 685600 110000 687000
rect 111600 685600 113000 687000
rect 114600 685600 116000 687000
rect 117600 685600 119000 687000
rect 120600 685600 122000 687000
rect 123600 685600 125000 687000
rect 126600 685600 128000 687000
rect 129600 685600 131000 687000
rect 132600 685600 134000 687000
rect 135600 685600 137000 687000
rect 138600 685600 140000 687000
rect 141600 685600 143000 687000
rect 144600 685600 146000 687000
rect 147600 685600 149000 687000
rect 150600 685600 152000 687000
rect 153600 685600 155000 687000
rect 156600 685600 158000 687000
rect 159600 685600 161000 687000
rect 162600 685600 164000 687000
rect 165600 685600 167000 687000
rect 168600 685600 170000 687000
rect 171600 685600 173000 687000
rect 174600 685600 176000 687000
rect 177600 685600 179000 687000
rect 180600 685600 182000 687000
rect 183600 685600 185000 687000
rect 186600 685600 188000 687000
rect 189600 685600 191000 687000
rect 192600 685600 194000 687000
rect 195600 685600 197000 687000
rect 198600 685600 200000 687000
rect 201600 685600 203000 687000
rect 204600 685600 206000 687000
rect 207600 685600 209000 687000
rect 210600 685600 212000 687000
rect 213600 685600 215000 687000
rect 216600 685600 218000 687000
rect 219600 685600 221000 687000
rect 222600 685600 224000 687000
rect 225600 685600 227000 687000
rect 228600 685600 230000 687000
rect 231600 685600 233000 687000
rect 234600 685600 236000 687000
rect 237600 685600 239000 687000
rect 240600 685600 242000 687000
rect 243600 685600 245000 687000
rect 246600 685600 248000 687000
rect 249600 685600 251000 687000
rect 252600 685600 254000 687000
rect 255600 685600 257000 687000
rect 258600 685600 260000 687000
rect 261600 685600 263000 687000
rect 264600 685600 266000 687000
rect 267600 685600 269000 687000
rect 270600 685600 272000 687000
rect 273600 685600 275000 687000
rect 276600 685600 278000 687000
rect 279600 685600 281000 687000
rect 282600 685600 284000 687000
rect 285600 685600 287000 687000
rect 288600 685600 290000 687000
rect 291600 685600 293000 687000
rect 294600 685600 296000 687000
rect 297600 685600 299000 687000
rect 300600 685600 302000 687000
rect 303600 685600 305000 687000
rect 306600 685600 308000 687000
rect 309600 685600 311000 687000
rect 312600 685600 314000 687000
rect 315600 685600 317000 687000
rect 318600 685600 320000 687000
rect 321600 685600 323000 687000
rect 324600 685600 326000 687000
rect 327600 685600 329000 687000
rect 330600 685600 332000 687000
rect 333600 685600 335000 687000
rect 336600 685600 338000 687000
rect 339600 685600 341000 687000
rect 342600 685600 344000 687000
rect 345600 685600 347000 687000
rect 348600 685600 350000 687000
rect 351600 685600 353000 687000
rect 354600 685600 356000 687000
rect 357600 685600 359000 687000
rect 360600 685600 362000 687000
rect 363600 685600 365000 687000
rect 366600 685600 368000 687000
rect 369600 685600 371000 687000
rect 372600 685600 374000 687000
rect 375600 685600 377000 687000
rect 378600 685600 380000 687000
rect 381600 685600 383000 687000
rect 384600 685600 386000 687000
rect 387600 685600 389000 687000
rect 390600 685600 392000 687000
rect 393600 685600 395000 687000
rect 396600 685600 398000 687000
rect 399600 685600 401000 687000
rect 402600 685600 404000 687000
rect 405600 685600 407000 687000
rect 408600 685600 410000 687000
rect 411600 685600 413000 687000
rect 414600 685600 416000 687000
rect 417600 685600 419000 687000
rect 420600 685600 422000 687000
rect 423600 685600 425000 687000
rect 426600 685600 428000 687000
rect 429600 685600 431000 687000
rect 432600 685600 434000 687000
rect 435600 685600 437000 687000
rect 438600 685600 440000 687000
rect 441600 685600 443000 687000
rect 444600 685600 446000 687000
rect 447600 685600 449000 687000
rect 450600 685600 452000 687000
rect 453600 685600 455000 687000
rect 456600 685600 458000 687000
rect 459600 685600 461000 687000
rect 462600 685600 464000 687000
rect 465600 685600 467000 687000
rect 468600 685600 470000 687000
rect 471600 685600 473000 687000
rect 474600 685600 476000 687000
rect 477600 685600 479000 687000
rect 480600 685600 482000 687000
rect 483600 685600 485000 687000
rect 486600 685600 488000 687000
rect 489600 685600 491000 687000
rect 492600 685600 494000 687000
rect 495600 685600 497000 687000
rect 498600 685600 500000 687000
rect 501600 685600 503000 687000
rect 504600 685600 506000 687000
rect 507600 685600 509000 687000
rect 510600 685600 512000 687000
rect 513600 685600 515000 687000
rect 516600 685600 518000 687000
rect 519600 685600 521000 687000
rect 522600 685600 524000 687000
rect 525600 685600 526600 687000
rect 4400 684000 526600 685600
rect 4400 682600 5400 684000
rect 7000 682600 9200 684000
rect 10800 682600 14000 684000
rect 15600 682600 17000 684000
rect 18600 682600 20000 684000
rect 21600 682600 23000 684000
rect 24600 682600 26000 684000
rect 27600 682600 29000 684000
rect 30600 682600 32000 684000
rect 33600 682600 35000 684000
rect 36600 682600 38000 684000
rect 39600 682600 41000 684000
rect 42600 682600 44000 684000
rect 45600 682600 47000 684000
rect 48600 682600 50000 684000
rect 51600 682600 53000 684000
rect 54600 682600 56000 684000
rect 57600 682600 59000 684000
rect 60600 682600 62000 684000
rect 63600 682600 65000 684000
rect 66600 682600 68000 684000
rect 69600 682600 71000 684000
rect 72600 682600 74000 684000
rect 75600 682600 77000 684000
rect 78600 682600 80000 684000
rect 81600 682600 83000 684000
rect 84600 682600 86000 684000
rect 87600 682600 89000 684000
rect 90600 682600 92000 684000
rect 93600 682600 95000 684000
rect 96600 682600 98000 684000
rect 99600 682600 101000 684000
rect 102600 682600 104000 684000
rect 105600 682600 107000 684000
rect 108600 682600 110000 684000
rect 111600 682600 113000 684000
rect 114600 682600 116000 684000
rect 117600 682600 119000 684000
rect 120600 682600 122000 684000
rect 123600 682600 125000 684000
rect 126600 682600 128000 684000
rect 129600 682600 131000 684000
rect 132600 682600 134000 684000
rect 135600 682600 137000 684000
rect 138600 682600 140000 684000
rect 141600 682600 143000 684000
rect 144600 682600 146000 684000
rect 147600 682600 149000 684000
rect 150600 682600 152000 684000
rect 153600 682600 155000 684000
rect 156600 682600 158000 684000
rect 159600 682600 161000 684000
rect 162600 682600 164000 684000
rect 165600 682600 167000 684000
rect 168600 682600 170000 684000
rect 171600 682600 173000 684000
rect 174600 682600 176000 684000
rect 177600 682600 179000 684000
rect 180600 682600 182000 684000
rect 183600 682600 185000 684000
rect 186600 682600 188000 684000
rect 189600 682600 191000 684000
rect 192600 682600 194000 684000
rect 195600 682600 197000 684000
rect 198600 682600 200000 684000
rect 201600 682600 203000 684000
rect 204600 682600 206000 684000
rect 207600 682600 209000 684000
rect 210600 682600 212000 684000
rect 213600 682600 215000 684000
rect 216600 682600 218000 684000
rect 219600 682600 221000 684000
rect 222600 682600 224000 684000
rect 225600 682600 227000 684000
rect 228600 682600 230000 684000
rect 231600 682600 233000 684000
rect 234600 682600 236000 684000
rect 237600 682600 239000 684000
rect 240600 682600 242000 684000
rect 243600 682600 245000 684000
rect 246600 682600 248000 684000
rect 249600 682600 251000 684000
rect 252600 682600 254000 684000
rect 255600 682600 257000 684000
rect 258600 682600 260000 684000
rect 261600 682600 263000 684000
rect 264600 682600 266000 684000
rect 267600 682600 269000 684000
rect 270600 682600 272000 684000
rect 273600 682600 275000 684000
rect 276600 682600 278000 684000
rect 279600 682600 281000 684000
rect 282600 682600 284000 684000
rect 285600 682600 287000 684000
rect 288600 682600 290000 684000
rect 291600 682600 293000 684000
rect 294600 682600 296000 684000
rect 297600 682600 299000 684000
rect 300600 682600 302000 684000
rect 303600 682600 305000 684000
rect 306600 682600 308000 684000
rect 309600 682600 311000 684000
rect 312600 682600 314000 684000
rect 315600 682600 317000 684000
rect 318600 682600 320000 684000
rect 321600 682600 323000 684000
rect 324600 682600 326000 684000
rect 327600 682600 329000 684000
rect 330600 682600 332000 684000
rect 333600 682600 335000 684000
rect 336600 682600 338000 684000
rect 339600 682600 341000 684000
rect 342600 682600 344000 684000
rect 345600 682600 347000 684000
rect 348600 682600 350000 684000
rect 351600 682600 353000 684000
rect 354600 682600 356000 684000
rect 357600 682600 359000 684000
rect 360600 682600 362000 684000
rect 363600 682600 365000 684000
rect 366600 682600 368000 684000
rect 369600 682600 371000 684000
rect 372600 682600 374000 684000
rect 375600 682600 377000 684000
rect 378600 682600 380000 684000
rect 381600 682600 383000 684000
rect 384600 682600 386000 684000
rect 387600 682600 389000 684000
rect 390600 682600 392000 684000
rect 393600 682600 395000 684000
rect 396600 682600 398000 684000
rect 399600 682600 401000 684000
rect 402600 682600 404000 684000
rect 405600 682600 407000 684000
rect 408600 682600 410000 684000
rect 411600 682600 413000 684000
rect 414600 682600 416000 684000
rect 417600 682600 419000 684000
rect 420600 682600 422000 684000
rect 423600 682600 425000 684000
rect 426600 682600 428000 684000
rect 429600 682600 431000 684000
rect 432600 682600 434000 684000
rect 435600 682600 437000 684000
rect 438600 682600 440000 684000
rect 441600 682600 443000 684000
rect 444600 682600 446000 684000
rect 447600 682600 449000 684000
rect 450600 682600 452000 684000
rect 453600 682600 455000 684000
rect 456600 682600 458000 684000
rect 459600 682600 461000 684000
rect 462600 682600 464000 684000
rect 465600 682600 467000 684000
rect 468600 682600 470000 684000
rect 471600 682600 473000 684000
rect 474600 682600 476000 684000
rect 477600 682600 479000 684000
rect 480600 682600 482000 684000
rect 483600 682600 485000 684000
rect 486600 682600 488000 684000
rect 489600 682600 491000 684000
rect 492600 682600 494000 684000
rect 495600 682600 497000 684000
rect 498600 682600 500000 684000
rect 501600 682600 503000 684000
rect 504600 682600 506000 684000
rect 507600 682600 509000 684000
rect 510600 682600 512000 684000
rect 513600 682600 515000 684000
rect 516600 682600 518000 684000
rect 519600 682600 521000 684000
rect 522600 682600 524000 684000
rect 525600 682600 526600 684000
rect 4400 681000 526600 682600
rect 4400 679600 5400 681000
rect 7000 679600 9200 681000
rect 10800 679600 14000 681000
rect 15600 679600 526600 681000
rect 4400 678000 16600 679600
rect 4400 676600 5400 678000
rect 7000 676600 9200 678000
rect 10800 676600 14000 678000
rect 15600 676600 16600 678000
rect 510000 677400 526600 679600
rect 580110 682990 583580 683510
rect 580110 678030 580470 682990
rect 581910 678030 583580 682990
rect 580110 677660 583580 678030
rect 4400 675000 16600 676600
rect 4400 673600 5400 675000
rect 7000 673600 9200 675000
rect 10800 673600 14000 675000
rect 15600 673600 16600 675000
rect 4400 672000 16600 673600
rect 4400 670600 5400 672000
rect 7000 670600 9200 672000
rect 10800 670600 14000 672000
rect 15600 670600 16600 672000
rect 4400 669000 16600 670600
rect 4400 667600 5400 669000
rect 7000 667600 9200 669000
rect 10800 667600 14000 669000
rect 15600 667600 16600 669000
rect 519680 669740 527080 670340
rect 4400 666000 16600 667600
rect 498570 668160 514790 668240
rect 498570 668100 512660 668160
rect 498570 667090 498670 668100
rect 500420 667690 512660 668100
rect 513650 667690 514790 668160
rect 500420 667610 514790 667690
rect 500420 667090 500530 667610
rect 498570 666930 500530 667090
rect 514270 666530 514790 667610
rect 4400 664600 5400 666000
rect 7000 664600 9200 666000
rect 10800 664600 14000 666000
rect 15600 664600 16600 666000
rect 503960 665340 514800 665370
rect 4400 663000 16600 664600
rect 503850 665300 514800 665340
rect 503850 665220 514320 665300
rect 503850 664910 512420 665220
rect 514020 664910 514320 665220
rect 503850 664830 514320 664910
rect 514680 664830 514800 665300
rect 503850 664810 514800 664830
rect 503850 664210 504430 664810
rect 519680 664340 520580 669740
rect 526480 664340 527080 669740
rect 4400 661600 5400 663000
rect 7000 661600 9200 663000
rect 10800 661600 14000 663000
rect 15600 661600 16600 663000
rect 4400 660000 16600 661600
rect 503900 660260 504400 664210
rect 519680 663640 527080 664340
rect 4400 658600 5400 660000
rect 7000 658600 9200 660000
rect 10800 658600 14000 660000
rect 15600 658600 16600 660000
rect 4400 657000 16600 658600
rect 4400 655600 5400 657000
rect 7000 655600 9200 657000
rect 10800 655600 14000 657000
rect 15600 655600 16600 657000
rect 503880 658200 504400 660260
rect 4400 654000 16600 655600
rect 4400 652600 5400 654000
rect 7000 652600 9200 654000
rect 10800 652600 14000 654000
rect 15600 652600 16600 654000
rect 4400 651000 16600 652600
rect 499320 654350 499710 655980
rect 503880 654350 504380 658200
rect 505780 656570 511880 656640
rect 499320 653910 504380 654350
rect 505160 654640 511880 656570
rect 505160 654000 506330 654640
rect 499320 652230 499710 653910
rect 4400 649600 5400 651000
rect 7000 649600 9200 651000
rect 10800 649600 14000 651000
rect 15600 649600 16600 651000
rect 4400 648000 16600 649600
rect 4400 646600 5400 648000
rect 7000 646600 9200 648000
rect 10800 646600 14000 648000
rect 15600 646600 16600 648000
rect 4400 645000 16600 646600
rect 4400 643600 5400 645000
rect 7000 643600 9200 645000
rect 10800 643600 14000 645000
rect 15600 643600 16600 645000
rect 4400 642000 16600 643600
rect 4400 640600 5400 642000
rect 7000 640600 9200 642000
rect 10800 640600 14000 642000
rect 15600 640600 16600 642000
rect 4400 639000 16600 640600
rect 4400 637600 5400 639000
rect 7000 637600 9200 639000
rect 10800 637600 14000 639000
rect 15600 637600 16600 639000
rect 4400 636000 16600 637600
rect 4400 634600 5400 636000
rect 7000 634600 9200 636000
rect 10800 634600 14000 636000
rect 15600 634600 16600 636000
rect 4400 633000 16600 634600
rect 4400 631600 5400 633000
rect 7000 631600 9200 633000
rect 10800 631600 14000 633000
rect 15600 631600 16600 633000
rect 4400 630000 16600 631600
rect 4400 628600 5400 630000
rect 7000 628600 9200 630000
rect 10800 628600 14000 630000
rect 15600 628600 16600 630000
rect 4400 627000 16600 628600
rect 4400 625600 5400 627000
rect 7000 625600 9200 627000
rect 10800 625600 14000 627000
rect 15600 625600 16600 627000
rect 4400 624000 16600 625600
rect 4400 622600 5400 624000
rect 7000 622600 9200 624000
rect 10800 622600 14000 624000
rect 15600 622600 16600 624000
rect 4400 621000 16600 622600
rect 4400 619600 5400 621000
rect 7000 619600 9200 621000
rect 10800 619600 14000 621000
rect 15600 619600 16600 621000
rect 4400 618000 16600 619600
rect 4400 616600 5400 618000
rect 7000 616600 9200 618000
rect 10800 616600 14000 618000
rect 15600 616600 16600 618000
rect 509180 623740 511880 654640
rect 519780 646740 527180 647440
rect 519780 641340 520780 646740
rect 526680 641340 527180 646740
rect 519780 640740 527180 641340
rect 576350 644270 583900 644590
rect 576350 630020 576690 644270
rect 583530 630020 583900 644270
rect 576350 629740 583900 630020
rect 509180 623040 527180 623740
rect 509180 617740 520580 623040
rect 526580 617740 527180 623040
rect 509180 617040 527180 617740
rect 4400 615000 16600 616600
rect 4400 613600 5400 615000
rect 7000 613600 9200 615000
rect 10800 613600 14000 615000
rect 15600 613600 16600 615000
rect 4400 612000 16600 613600
rect 4400 610600 5400 612000
rect 7000 610600 9200 612000
rect 10800 610600 14000 612000
rect 15600 610600 16600 612000
rect 4400 609000 16600 610600
rect 4400 607600 5400 609000
rect 7000 607600 9200 609000
rect 10800 607600 14000 609000
rect 15600 607600 16600 609000
rect 4400 606000 16600 607600
rect 4400 604600 5400 606000
rect 7000 604600 9200 606000
rect 10800 604600 14000 606000
rect 15600 604600 16600 606000
rect 4400 603000 16600 604600
rect 4400 601600 5400 603000
rect 7000 601600 9200 603000
rect 10800 601600 14000 603000
rect 15600 601600 16600 603000
rect 4400 600000 16600 601600
rect 4400 598600 5400 600000
rect 7000 598600 9200 600000
rect 10800 598600 14000 600000
rect 15600 598600 16600 600000
rect 4400 597000 16600 598600
rect 4400 595600 5400 597000
rect 7000 595600 9200 597000
rect 10800 595600 14000 597000
rect 15600 595600 16600 597000
rect 4400 594000 16600 595600
rect 4400 592600 5400 594000
rect 7000 592600 9200 594000
rect 10800 592600 14000 594000
rect 15600 592600 16600 594000
rect 4400 591000 16600 592600
rect 4400 589600 5400 591000
rect 7000 589600 9200 591000
rect 10800 589600 14000 591000
rect 15600 589600 16600 591000
rect 4400 588000 16600 589600
rect 4400 586600 5400 588000
rect 7000 586600 9200 588000
rect 10800 586600 14000 588000
rect 15600 586600 16600 588000
rect 4400 585000 16600 586600
rect 4400 583600 5400 585000
rect 7000 583600 9200 585000
rect 10800 583600 14000 585000
rect 15600 583600 16600 585000
rect 4400 582000 16600 583600
rect 4400 580600 5400 582000
rect 7000 580600 9200 582000
rect 10800 580600 14000 582000
rect 15600 580600 16600 582000
rect 4400 579000 16600 580600
rect 577270 583570 583810 584240
rect 577270 580390 577730 583570
rect 583180 580390 583810 583570
rect 577270 579860 583810 580390
rect 4400 577600 5400 579000
rect 7000 577600 9200 579000
rect 10800 577600 14000 579000
rect 15600 577600 16600 579000
rect 4400 576000 16600 577600
rect 4400 574600 5400 576000
rect 7000 574600 9200 576000
rect 10800 574600 14000 576000
rect 15600 574600 16600 576000
rect 4400 573000 16600 574600
rect 4400 571600 5400 573000
rect 7000 571600 9200 573000
rect 10800 571600 14000 573000
rect 15600 571600 16600 573000
rect 511690 574080 519090 574680
rect 4400 570000 16600 571600
rect 490580 572500 507000 572580
rect 490580 572440 504870 572500
rect 490580 571430 490680 572440
rect 492430 572030 504870 572440
rect 505860 572030 507000 572500
rect 492430 571950 507000 572030
rect 492430 571430 492540 571950
rect 490580 571270 492540 571430
rect 506480 570870 507000 571950
rect 4400 568600 5400 570000
rect 7000 568600 9200 570000
rect 10800 568600 14000 570000
rect 15600 568600 16600 570000
rect 495970 569680 507010 569710
rect 4400 567000 16600 568600
rect 495860 569640 507010 569680
rect 495860 569560 506530 569640
rect 495860 569250 504630 569560
rect 506230 569250 506530 569560
rect 495860 569170 506530 569250
rect 506890 569170 507010 569640
rect 495860 569150 507010 569170
rect 495860 568550 496440 569150
rect 511690 568680 512590 574080
rect 518490 568680 519090 574080
rect 564280 574210 571680 574810
rect 543170 572630 559590 572710
rect 543170 572570 557460 572630
rect 543170 571560 543270 572570
rect 545020 572160 557460 572570
rect 558450 572160 559590 572630
rect 545020 572080 559590 572160
rect 545020 571560 545130 572080
rect 543170 571400 545130 571560
rect 548560 569810 559600 569840
rect 548450 569770 559600 569810
rect 548450 569690 559120 569770
rect 548450 569380 557220 569690
rect 558820 569380 559120 569690
rect 548450 569300 559120 569380
rect 559480 569300 559600 569770
rect 548450 569280 559600 569300
rect 548450 568680 549030 569280
rect 564280 568810 565180 574210
rect 571080 568810 571680 574210
rect 4400 565600 5400 567000
rect 7000 565600 9200 567000
rect 10800 565600 14000 567000
rect 15600 565600 16600 567000
rect 4400 564800 16600 565600
rect 1200 564730 17600 564800
rect 330 564400 17600 564730
rect 495910 564600 496410 568550
rect 511690 567980 519090 568680
rect 548500 564730 549000 568680
rect 564280 568110 571680 568810
rect 330 564320 4400 564400
rect 330 549250 870 564320
rect 2600 563000 4400 564320
rect 6000 563000 7200 564400
rect 8800 563000 9800 564400
rect 11400 563000 12800 564400
rect 14400 563000 15600 564400
rect 17200 563000 17600 564400
rect 2600 561400 17600 563000
rect 2600 560000 4400 561400
rect 6000 560000 7200 561400
rect 8800 560000 9800 561400
rect 11400 560000 12800 561400
rect 14400 560000 15600 561400
rect 17200 560000 17600 561400
rect 495890 562540 496410 564600
rect 548480 562670 549000 564730
rect 2600 558200 17600 560000
rect 2600 556800 4400 558200
rect 6000 556800 7200 558200
rect 8800 556800 9800 558200
rect 11400 556800 12800 558200
rect 14400 556800 15600 558200
rect 17200 556800 17600 558200
rect 2600 555800 17600 556800
rect 491330 558690 491720 560320
rect 495890 558690 496390 562540
rect 497790 560910 503890 560980
rect 491330 558250 496390 558690
rect 497170 558980 503890 560910
rect 497170 558340 498340 558980
rect 491330 556570 491720 558250
rect 2600 554400 4400 555800
rect 6000 554400 7200 555800
rect 8800 554400 9800 555800
rect 11400 554400 12800 555800
rect 14400 554400 15600 555800
rect 17200 554400 17600 555800
rect 2600 553200 17600 554400
rect 2600 551800 4400 553200
rect 6000 551800 7200 553200
rect 8800 551800 9800 553200
rect 11400 551800 12800 553200
rect 14400 551800 15600 553200
rect 17200 551800 17600 553200
rect 2600 551600 16000 551800
rect 16600 551600 17600 551800
rect 2600 550600 17600 551600
rect 2600 549250 4400 550600
rect 330 549200 4400 549250
rect 6000 549200 7200 550600
rect 8800 549200 9800 550600
rect 11400 549200 12800 550600
rect 14400 549200 15600 550600
rect 17200 549200 17600 550600
rect 330 548720 16000 549200
rect 1200 548600 16000 548720
rect 16600 548600 17600 549200
rect 1200 548400 17600 548600
rect 6880 536700 7340 536740
rect 6880 534720 6920 536700
rect 7200 534720 7340 536700
rect 6880 534680 7340 534720
rect 8380 536700 8740 536740
rect 8380 534720 8420 536700
rect 8700 534720 8740 536700
rect 8380 534680 8740 534720
rect 501190 528080 503890 558980
rect 543920 558820 544310 560450
rect 548480 558820 548980 562670
rect 550380 561040 556480 561110
rect 543920 558380 548980 558820
rect 549760 559110 556480 561040
rect 549760 558470 550930 559110
rect 543920 556700 544310 558380
rect 511790 551080 519190 551780
rect 511790 545680 512790 551080
rect 518690 545680 519190 551080
rect 511790 545080 519190 545680
rect 553780 528210 556480 559110
rect 564380 551210 571780 551910
rect 564380 545810 565380 551210
rect 571280 545810 571780 551210
rect 564380 545210 571780 545810
rect 501190 527380 519190 528080
rect 501190 522080 512590 527380
rect 518590 522080 519190 527380
rect 501190 521380 519190 522080
rect 553780 527510 571780 528210
rect 553780 522210 565180 527510
rect 571180 522210 571780 527510
rect 553780 521510 571780 522210
rect 160 512460 2530 512620
rect 160 511100 300 512460
rect 2350 511100 2530 512460
rect 160 510950 2530 511100
rect 567980 501420 569290 501520
rect 553280 500380 557030 500770
rect 554960 496210 555400 500380
rect 567980 499670 568140 501420
rect 569150 499670 569290 501420
rect 567980 499560 569290 499670
rect 554960 496190 561310 496210
rect 565260 496190 566390 496240
rect 554960 496130 566390 496190
rect 554960 495710 566420 496130
rect 559250 495690 566420 495710
rect 565260 495660 566420 495690
rect 555050 494310 557620 494930
rect 555050 493760 557690 494310
rect 555690 490910 557690 493760
rect 518090 488210 557690 490910
rect 518090 479510 524790 488210
rect 565860 487470 566420 495660
rect 565860 485870 565960 487470
rect 566270 485870 566420 487470
rect 565860 485570 566420 485870
rect 565860 485210 565880 485570
rect 566350 485210 566420 485570
rect 565860 485090 566420 485210
rect 568660 487230 569290 499560
rect 580300 495690 582680 496130
rect 580300 493390 580590 495690
rect 582340 493390 582680 495690
rect 580300 493190 582680 493390
rect 568660 486240 568740 487230
rect 569210 486240 569290 487230
rect 568660 485100 569290 486240
rect 518090 473510 518790 479510
rect 524090 473510 524790 479510
rect 518090 472910 524790 473510
rect 541790 479310 548490 480310
rect 541790 473410 542390 479310
rect 547790 473410 548490 479310
rect 541790 472910 548490 473410
rect 564690 479510 571390 480410
rect 564690 473610 565390 479510
rect 570790 473610 571390 479510
rect 564690 473010 571390 473610
rect 190 469210 2560 469370
rect 190 467850 330 469210
rect 2380 467850 2560 469210
rect 190 467700 2560 467850
rect 576460 450970 578840 451410
rect 576460 448670 576750 450970
rect 578500 448670 578840 450970
rect 576460 448470 578840 448670
rect 200 424600 2000 424800
rect 200 423400 400 424600
rect 1800 423400 2000 424600
rect 200 423200 2000 423400
rect 571350 407140 583800 407350
rect 571350 405820 571720 407140
rect 577750 405820 583800 407140
rect 571350 405610 583800 405820
rect 200 381300 2200 381500
rect 200 380100 400 381300
rect 1800 380100 2200 381300
rect 200 379900 2200 380100
rect 900 370900 2200 379900
rect 300 369000 2200 370900
rect 300 342310 1500 369000
rect 575600 365000 576200 365200
rect 578400 365000 579000 365200
rect 573800 364800 574800 365000
rect 573800 363400 574000 364800
rect 574600 363400 574800 364800
rect 573800 363200 574800 363400
rect 575600 363400 575800 365000
rect 576000 363400 576200 365000
rect 575600 363200 576200 363400
rect 576600 364800 577600 365000
rect 576600 363400 576800 364800
rect 577400 363400 577600 364800
rect 576600 363200 577600 363400
rect 578400 363400 578600 365000
rect 578800 363400 579000 365000
rect 578400 363200 579000 363400
rect 572400 361400 574800 361800
rect 572400 361200 572600 361400
rect 573400 361200 573800 361400
rect 574600 361240 574800 361400
rect 574600 361200 575900 361240
rect 572400 361000 575900 361200
rect 572400 360800 572600 361000
rect 573400 360800 573800 361000
rect 574600 360800 575900 361000
rect 572400 360600 575900 360800
rect 572400 360400 572600 360600
rect 573400 360400 573800 360600
rect 574600 360400 575900 360600
rect 572400 360200 575900 360400
rect 572400 360000 572600 360200
rect 573400 360000 573800 360200
rect 574600 360000 575900 360200
rect 572400 359800 575900 360000
rect 572400 359600 572600 359800
rect 573400 359600 573800 359800
rect 574600 359600 575900 359800
rect 572400 359400 575900 359600
rect 572400 359200 572600 359400
rect 573400 359200 573800 359400
rect 574600 359200 575900 359400
rect 579020 360800 583790 360900
rect 579020 359440 579150 360800
rect 582190 359440 583790 360800
rect 579020 359300 583790 359440
rect 572400 359000 575900 359200
rect 572400 358800 572600 359000
rect 573400 358800 573800 359000
rect 574600 358800 575900 359000
rect 572400 358600 575900 358800
rect 572400 358400 572600 358600
rect 573400 358400 573800 358600
rect 574600 358400 575900 358600
rect 572400 358200 575900 358400
rect 572400 358000 572600 358200
rect 573400 358000 573800 358200
rect 574600 358000 575900 358200
rect 572400 357800 575900 358000
rect 572400 357600 572600 357800
rect 573400 357600 573800 357800
rect 574600 357600 575900 357800
rect 572400 357400 575900 357600
rect 572400 357200 572600 357400
rect 573400 357200 573800 357400
rect 574600 357200 575900 357400
rect 572400 357000 575900 357200
rect 572400 356800 572600 357000
rect 573400 356800 573800 357000
rect 574600 356800 575900 357000
rect 572400 356600 575900 356800
rect 572400 356400 572600 356600
rect 573400 356400 573800 356600
rect 574600 356400 575900 356600
rect 572400 356200 575900 356400
rect 572400 356000 572600 356200
rect 573400 356000 573800 356200
rect 574600 356000 575900 356200
rect 572400 355800 575900 356000
rect 572400 355600 572600 355800
rect 573400 355600 573800 355800
rect 574600 355600 575900 355800
rect 572400 355400 575900 355600
rect 572400 355200 572600 355400
rect 573400 355200 573800 355400
rect 574600 355200 575900 355400
rect 572400 355000 575900 355200
rect 572400 354800 572600 355000
rect 573400 354800 573800 355000
rect 574600 354800 575900 355000
rect 572400 354760 575900 354800
rect 572400 354600 574800 354760
rect 572400 354400 572600 354600
rect 573400 354400 573800 354600
rect 574600 354400 574800 354600
rect 572400 354200 574800 354400
rect 572400 354000 572600 354200
rect 573400 354000 573800 354200
rect 574600 354000 574800 354200
rect 572400 353800 574800 354000
rect 576020 354520 576520 354560
rect 576020 354460 576050 354520
rect 576180 354460 576520 354520
rect 576020 353350 576520 354460
rect 10083 343040 10473 344720
rect 3463 342310 4633 342950
rect 300 340400 4633 342310
rect 4500 340380 4633 340400
rect 5413 342600 10473 343040
rect 5413 338750 5913 342600
rect 10083 340970 10473 342600
rect 200 338100 2000 338300
rect 200 336900 400 338100
rect 1800 336900 2000 338100
rect 200 336700 2000 336900
rect 5393 336690 5913 338750
rect 5393 332740 5893 336690
rect 5363 332140 5943 332740
rect 2790 331610 5943 332140
rect 2790 331580 5833 331610
rect 2830 327510 3420 331580
rect 9270 330020 11240 330040
rect 9263 329860 11240 330020
rect 9263 329630 9373 329860
rect 9263 329340 9360 329630
rect 9260 328710 9360 329340
rect 11123 328850 11240 329860
rect 2830 326413 3390 327510
rect 9270 327350 9360 328710
rect 2830 324813 2930 326413
rect 3240 324813 3390 326413
rect 2830 324513 3390 324813
rect 2830 324153 2850 324513
rect 3320 324153 3390 324513
rect 2830 324033 3390 324153
rect 5630 326173 9360 327350
rect 5630 325183 5710 326173
rect 6180 325183 9360 326173
rect 5630 324140 9360 325183
rect 5630 324043 6260 324140
rect 9270 324110 9360 324140
rect 11100 324110 11240 328850
rect 9270 323850 11240 324110
rect 3600 323000 8500 323200
rect 3600 322000 3800 323000
rect 7400 322000 8500 323000
rect 3600 321800 8500 322000
rect 200 296100 2000 296300
rect 200 294900 400 296100
rect 1800 294900 2000 296100
rect 200 294700 2000 294900
rect 200 253000 2000 253200
rect 200 251800 400 253000
rect 1800 251800 2000 253000
rect 200 251600 2000 251800
rect 400 177370 2740 177720
rect 400 163110 700 177370
rect 2330 163110 2740 177370
rect 400 162870 2740 163110
rect 6100 125700 8500 321800
rect 573520 271200 576520 353350
rect 576860 354530 577330 354570
rect 576860 354450 577180 354530
rect 577310 354450 577330 354530
rect 576860 353350 577330 354450
rect 576860 315640 579860 353350
rect 576850 315490 583800 315640
rect 576850 314100 576980 315490
rect 579620 314100 583800 315490
rect 576850 313990 583800 314100
rect 576860 312370 579860 313990
rect 573510 270990 583830 271200
rect 573510 269790 573690 270990
rect 579290 269790 583830 270990
rect 573510 269620 583830 269790
rect 573520 269100 576520 269620
rect 576000 215950 576390 217650
rect 569160 215220 571600 215910
rect 576000 215600 577440 215950
rect 569150 131380 571600 215220
rect 577050 213900 577440 215600
rect 579200 201000 581200 201200
rect 579200 198160 579460 201000
rect 580960 198160 581200 201000
rect 579200 189900 579500 198160
rect 580900 189900 581200 198160
rect 579200 189500 581200 189900
rect 576200 175500 579600 175800
rect 576200 167200 576400 175500
rect 579400 167200 579600 175500
rect 576200 166600 579600 167200
rect 572900 152000 576700 152600
rect 572900 151830 573200 152000
rect 572900 148990 573150 151830
rect 572900 143700 573200 148990
rect 576200 143700 576700 152000
rect 572900 143300 576700 143700
rect 569150 131300 575820 131380
rect 569150 130820 577940 131300
rect 569150 130770 570880 130820
rect 569150 128110 570850 130770
rect 200 125500 8500 125700
rect 200 124300 400 125500
rect 1800 124300 8500 125500
rect 200 124100 8500 124300
rect 569270 123400 570850 128110
rect 577350 123400 577940 130820
rect 569270 122970 577940 123400
rect 571390 122890 577940 122970
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 15690 701230 21540 703180
rect 67850 701700 73380 703110
rect 228670 701850 232530 702520
rect 330480 701740 334340 702410
rect 463720 699400 471140 701590
rect 510880 696600 525130 703440
rect 566440 699450 573030 701120
rect 5400 691600 7000 693000
rect 9200 691600 10800 693000
rect 14000 691600 15600 693000
rect 17000 691600 18600 693000
rect 20000 691600 21600 693000
rect 23000 691600 24600 693000
rect 26000 691600 27600 693000
rect 29000 691600 30600 693000
rect 32000 691600 33600 693000
rect 35000 691600 36600 693000
rect 38000 691600 39600 693000
rect 41000 691600 42600 693000
rect 44000 691600 45600 693000
rect 47000 691600 48600 693000
rect 50000 691600 51600 693000
rect 53000 691600 54600 693000
rect 56000 691600 57600 693000
rect 59000 691600 60600 693000
rect 62000 691600 63600 693000
rect 65000 691600 66600 693000
rect 68000 691600 69600 693000
rect 71000 691600 72600 693000
rect 74000 691600 75600 693000
rect 77000 691600 78600 693000
rect 80000 691600 81600 693000
rect 83000 691600 84600 693000
rect 86000 691600 87600 693000
rect 89000 691600 90600 693000
rect 92000 691600 93600 693000
rect 95000 691600 96600 693000
rect 98000 691600 99600 693000
rect 101000 691600 102600 693000
rect 104000 691600 105600 693000
rect 107000 691600 108600 693000
rect 110000 691600 111600 693000
rect 113000 691600 114600 693000
rect 116000 691600 117600 693000
rect 119000 691600 120600 693000
rect 122000 691600 123600 693000
rect 125000 691600 126600 693000
rect 128000 691600 129600 693000
rect 131000 691600 132600 693000
rect 134000 691600 135600 693000
rect 137000 691600 138600 693000
rect 140000 691600 141600 693000
rect 143000 691600 144600 693000
rect 146000 691600 147600 693000
rect 149000 691600 150600 693000
rect 152000 691600 153600 693000
rect 155000 691600 156600 693000
rect 158000 691600 159600 693000
rect 161000 691600 162600 693000
rect 164000 691600 165600 693000
rect 167000 691600 168600 693000
rect 170000 691600 171600 693000
rect 173000 691600 174600 693000
rect 176000 691600 177600 693000
rect 179000 691600 180600 693000
rect 182000 691600 183600 693000
rect 185000 691600 186600 693000
rect 188000 691600 189600 693000
rect 191000 691600 192600 693000
rect 194000 691600 195600 693000
rect 197000 691600 198600 693000
rect 200000 691600 201600 693000
rect 203000 691600 204600 693000
rect 206000 691600 207600 693000
rect 209000 691600 210600 693000
rect 212000 691600 213600 693000
rect 215000 691600 216600 693000
rect 218000 691600 219600 693000
rect 221000 691600 222600 693000
rect 224000 691600 225600 693000
rect 227000 691600 228600 693000
rect 230000 691600 231600 693000
rect 233000 691600 234600 693000
rect 236000 691600 237600 693000
rect 239000 691600 240600 693000
rect 242000 691600 243600 693000
rect 245000 691600 246600 693000
rect 248000 691600 249600 693000
rect 251000 691600 252600 693000
rect 254000 691600 255600 693000
rect 257000 691600 258600 693000
rect 260000 691600 261600 693000
rect 263000 691600 264600 693000
rect 266000 691600 267600 693000
rect 269000 691600 270600 693000
rect 272000 691600 273600 693000
rect 275000 691600 276600 693000
rect 278000 691600 279600 693000
rect 281000 691600 282600 693000
rect 284000 691600 285600 693000
rect 287000 691600 288600 693000
rect 290000 691600 291600 693000
rect 293000 691600 294600 693000
rect 296000 691600 297600 693000
rect 299000 691600 300600 693000
rect 302000 691600 303600 693000
rect 305000 691600 306600 693000
rect 308000 691600 309600 693000
rect 311000 691600 312600 693000
rect 314000 691600 315600 693000
rect 317000 691600 318600 693000
rect 320000 691600 321600 693000
rect 323000 691600 324600 693000
rect 326000 691600 327600 693000
rect 329000 691600 330600 693000
rect 332000 691600 333600 693000
rect 335000 691600 336600 693000
rect 338000 691600 339600 693000
rect 341000 691600 342600 693000
rect 344000 691600 345600 693000
rect 347000 691600 348600 693000
rect 350000 691600 351600 693000
rect 353000 691600 354600 693000
rect 356000 691600 357600 693000
rect 359000 691600 360600 693000
rect 362000 691600 363600 693000
rect 365000 691600 366600 693000
rect 368000 691600 369600 693000
rect 371000 691600 372600 693000
rect 374000 691600 375600 693000
rect 377000 691600 378600 693000
rect 380000 691600 381600 693000
rect 383000 691600 384600 693000
rect 386000 691600 387600 693000
rect 389000 691600 390600 693000
rect 392000 691600 393600 693000
rect 395000 691600 396600 693000
rect 398000 691600 399600 693000
rect 401000 691600 402600 693000
rect 404000 691600 405600 693000
rect 407000 691600 408600 693000
rect 410000 691600 411600 693000
rect 413000 691600 414600 693000
rect 416000 691600 417600 693000
rect 419000 691600 420600 693000
rect 422000 691600 423600 693000
rect 425000 691600 426600 693000
rect 428000 691600 429600 693000
rect 431000 691600 432600 693000
rect 434000 691600 435600 693000
rect 437000 691600 438600 693000
rect 440000 691600 441600 693000
rect 443000 691600 444600 693000
rect 446000 691600 447600 693000
rect 449000 691600 450600 693000
rect 452000 691600 453600 693000
rect 455000 691600 456600 693000
rect 458000 691600 459600 693000
rect 461000 691600 462600 693000
rect 464000 691600 465600 693000
rect 467000 691600 468600 693000
rect 470000 691600 471600 693000
rect 473000 691600 474600 693000
rect 476000 691600 477600 693000
rect 479000 691600 480600 693000
rect 482000 691600 483600 693000
rect 485000 691600 486600 693000
rect 488000 691600 489600 693000
rect 491000 691600 492600 693000
rect 494000 691600 495600 693000
rect 497000 691600 498600 693000
rect 500000 691600 501600 693000
rect 503000 691600 504600 693000
rect 506000 691600 507600 693000
rect 509000 691600 510600 693000
rect 512000 691600 513600 693000
rect 515000 691600 516600 693000
rect 518000 691600 519600 693000
rect 521000 691600 522600 693000
rect 524000 691600 525600 693000
rect 5400 688600 7000 690000
rect 9200 688600 10800 690000
rect 14000 688600 15600 690000
rect 17000 688600 18600 690000
rect 20000 688600 21600 690000
rect 23000 688600 24600 690000
rect 26000 688600 27600 690000
rect 29000 688600 30600 690000
rect 32000 688600 33600 690000
rect 35000 688600 36600 690000
rect 38000 688600 39600 690000
rect 41000 688600 42600 690000
rect 44000 688600 45600 690000
rect 47000 688600 48600 690000
rect 50000 688600 51600 690000
rect 53000 688600 54600 690000
rect 56000 688600 57600 690000
rect 59000 688600 60600 690000
rect 62000 688600 63600 690000
rect 65000 688600 66600 690000
rect 68000 688600 69600 690000
rect 71000 688600 72600 690000
rect 74000 688600 75600 690000
rect 77000 688600 78600 690000
rect 80000 688600 81600 690000
rect 83000 688600 84600 690000
rect 86000 688600 87600 690000
rect 89000 688600 90600 690000
rect 92000 688600 93600 690000
rect 95000 688600 96600 690000
rect 98000 688600 99600 690000
rect 101000 688600 102600 690000
rect 104000 688600 105600 690000
rect 107000 688600 108600 690000
rect 110000 688600 111600 690000
rect 113000 688600 114600 690000
rect 116000 688600 117600 690000
rect 119000 688600 120600 690000
rect 122000 688600 123600 690000
rect 125000 688600 126600 690000
rect 128000 688600 129600 690000
rect 131000 688600 132600 690000
rect 134000 688600 135600 690000
rect 137000 688600 138600 690000
rect 140000 688600 141600 690000
rect 143000 688600 144600 690000
rect 146000 688600 147600 690000
rect 149000 688600 150600 690000
rect 152000 688600 153600 690000
rect 155000 688600 156600 690000
rect 158000 688600 159600 690000
rect 161000 688600 162600 690000
rect 164000 688600 165600 690000
rect 167000 688600 168600 690000
rect 170000 688600 171600 690000
rect 173000 688600 174600 690000
rect 176000 688600 177600 690000
rect 179000 688600 180600 690000
rect 182000 688600 183600 690000
rect 185000 688600 186600 690000
rect 188000 688600 189600 690000
rect 191000 688600 192600 690000
rect 194000 688600 195600 690000
rect 197000 688600 198600 690000
rect 200000 688600 201600 690000
rect 203000 688600 204600 690000
rect 206000 688600 207600 690000
rect 209000 688600 210600 690000
rect 212000 688600 213600 690000
rect 215000 688600 216600 690000
rect 218000 688600 219600 690000
rect 221000 688600 222600 690000
rect 224000 688600 225600 690000
rect 227000 688600 228600 690000
rect 230000 688600 231600 690000
rect 233000 688600 234600 690000
rect 236000 688600 237600 690000
rect 239000 688600 240600 690000
rect 242000 688600 243600 690000
rect 245000 688600 246600 690000
rect 248000 688600 249600 690000
rect 251000 688600 252600 690000
rect 254000 688600 255600 690000
rect 257000 688600 258600 690000
rect 260000 688600 261600 690000
rect 263000 688600 264600 690000
rect 266000 688600 267600 690000
rect 269000 688600 270600 690000
rect 272000 688600 273600 690000
rect 275000 688600 276600 690000
rect 278000 688600 279600 690000
rect 281000 688600 282600 690000
rect 284000 688600 285600 690000
rect 287000 688600 288600 690000
rect 290000 688600 291600 690000
rect 293000 688600 294600 690000
rect 296000 688600 297600 690000
rect 299000 688600 300600 690000
rect 302000 688600 303600 690000
rect 305000 688600 306600 690000
rect 308000 688600 309600 690000
rect 311000 688600 312600 690000
rect 314000 688600 315600 690000
rect 317000 688600 318600 690000
rect 320000 688600 321600 690000
rect 323000 688600 324600 690000
rect 326000 688600 327600 690000
rect 329000 688600 330600 690000
rect 332000 688600 333600 690000
rect 335000 688600 336600 690000
rect 338000 688600 339600 690000
rect 341000 688600 342600 690000
rect 344000 688600 345600 690000
rect 347000 688600 348600 690000
rect 350000 688600 351600 690000
rect 353000 688600 354600 690000
rect 356000 688600 357600 690000
rect 359000 688600 360600 690000
rect 362000 688600 363600 690000
rect 365000 688600 366600 690000
rect 368000 688600 369600 690000
rect 371000 688600 372600 690000
rect 374000 688600 375600 690000
rect 377000 688600 378600 690000
rect 380000 688600 381600 690000
rect 383000 688600 384600 690000
rect 386000 688600 387600 690000
rect 389000 688600 390600 690000
rect 392000 688600 393600 690000
rect 395000 688600 396600 690000
rect 398000 688600 399600 690000
rect 401000 688600 402600 690000
rect 404000 688600 405600 690000
rect 407000 688600 408600 690000
rect 410000 688600 411600 690000
rect 413000 688600 414600 690000
rect 416000 688600 417600 690000
rect 419000 688600 420600 690000
rect 422000 688600 423600 690000
rect 425000 688600 426600 690000
rect 428000 688600 429600 690000
rect 431000 688600 432600 690000
rect 434000 688600 435600 690000
rect 437000 688600 438600 690000
rect 440000 688600 441600 690000
rect 443000 688600 444600 690000
rect 446000 688600 447600 690000
rect 449000 688600 450600 690000
rect 452000 688600 453600 690000
rect 455000 688600 456600 690000
rect 458000 688600 459600 690000
rect 461000 688600 462600 690000
rect 464000 688600 465600 690000
rect 467000 688600 468600 690000
rect 470000 688600 471600 690000
rect 473000 688600 474600 690000
rect 476000 688600 477600 690000
rect 479000 688600 480600 690000
rect 482000 688600 483600 690000
rect 485000 688600 486600 690000
rect 488000 688600 489600 690000
rect 491000 688600 492600 690000
rect 494000 688600 495600 690000
rect 497000 688600 498600 690000
rect 500000 688600 501600 690000
rect 503000 688600 504600 690000
rect 506000 688600 507600 690000
rect 509000 688600 510600 690000
rect 512000 688600 513600 690000
rect 515000 688600 516600 690000
rect 518000 688600 519600 690000
rect 521000 688600 522600 690000
rect 524000 688600 525600 690000
rect 1340 679860 3090 685550
rect 5400 685600 7000 687000
rect 9200 685600 10800 687000
rect 14000 685600 15600 687000
rect 17000 685600 18600 687000
rect 20000 685600 21600 687000
rect 23000 685600 24600 687000
rect 26000 685600 27600 687000
rect 29000 685600 30600 687000
rect 32000 685600 33600 687000
rect 35000 685600 36600 687000
rect 38000 685600 39600 687000
rect 41000 685600 42600 687000
rect 44000 685600 45600 687000
rect 47000 685600 48600 687000
rect 50000 685600 51600 687000
rect 53000 685600 54600 687000
rect 56000 685600 57600 687000
rect 59000 685600 60600 687000
rect 62000 685600 63600 687000
rect 65000 685600 66600 687000
rect 68000 685600 69600 687000
rect 71000 685600 72600 687000
rect 74000 685600 75600 687000
rect 77000 685600 78600 687000
rect 80000 685600 81600 687000
rect 83000 685600 84600 687000
rect 86000 685600 87600 687000
rect 89000 685600 90600 687000
rect 92000 685600 93600 687000
rect 95000 685600 96600 687000
rect 98000 685600 99600 687000
rect 101000 685600 102600 687000
rect 104000 685600 105600 687000
rect 107000 685600 108600 687000
rect 110000 685600 111600 687000
rect 113000 685600 114600 687000
rect 116000 685600 117600 687000
rect 119000 685600 120600 687000
rect 122000 685600 123600 687000
rect 125000 685600 126600 687000
rect 128000 685600 129600 687000
rect 131000 685600 132600 687000
rect 134000 685600 135600 687000
rect 137000 685600 138600 687000
rect 140000 685600 141600 687000
rect 143000 685600 144600 687000
rect 146000 685600 147600 687000
rect 149000 685600 150600 687000
rect 152000 685600 153600 687000
rect 155000 685600 156600 687000
rect 158000 685600 159600 687000
rect 161000 685600 162600 687000
rect 164000 685600 165600 687000
rect 167000 685600 168600 687000
rect 170000 685600 171600 687000
rect 173000 685600 174600 687000
rect 176000 685600 177600 687000
rect 179000 685600 180600 687000
rect 182000 685600 183600 687000
rect 185000 685600 186600 687000
rect 188000 685600 189600 687000
rect 191000 685600 192600 687000
rect 194000 685600 195600 687000
rect 197000 685600 198600 687000
rect 200000 685600 201600 687000
rect 203000 685600 204600 687000
rect 206000 685600 207600 687000
rect 209000 685600 210600 687000
rect 212000 685600 213600 687000
rect 215000 685600 216600 687000
rect 218000 685600 219600 687000
rect 221000 685600 222600 687000
rect 224000 685600 225600 687000
rect 227000 685600 228600 687000
rect 230000 685600 231600 687000
rect 233000 685600 234600 687000
rect 236000 685600 237600 687000
rect 239000 685600 240600 687000
rect 242000 685600 243600 687000
rect 245000 685600 246600 687000
rect 248000 685600 249600 687000
rect 251000 685600 252600 687000
rect 254000 685600 255600 687000
rect 257000 685600 258600 687000
rect 260000 685600 261600 687000
rect 263000 685600 264600 687000
rect 266000 685600 267600 687000
rect 269000 685600 270600 687000
rect 272000 685600 273600 687000
rect 275000 685600 276600 687000
rect 278000 685600 279600 687000
rect 281000 685600 282600 687000
rect 284000 685600 285600 687000
rect 287000 685600 288600 687000
rect 290000 685600 291600 687000
rect 293000 685600 294600 687000
rect 296000 685600 297600 687000
rect 299000 685600 300600 687000
rect 302000 685600 303600 687000
rect 305000 685600 306600 687000
rect 308000 685600 309600 687000
rect 311000 685600 312600 687000
rect 314000 685600 315600 687000
rect 317000 685600 318600 687000
rect 320000 685600 321600 687000
rect 323000 685600 324600 687000
rect 326000 685600 327600 687000
rect 329000 685600 330600 687000
rect 332000 685600 333600 687000
rect 335000 685600 336600 687000
rect 338000 685600 339600 687000
rect 341000 685600 342600 687000
rect 344000 685600 345600 687000
rect 347000 685600 348600 687000
rect 350000 685600 351600 687000
rect 353000 685600 354600 687000
rect 356000 685600 357600 687000
rect 359000 685600 360600 687000
rect 362000 685600 363600 687000
rect 365000 685600 366600 687000
rect 368000 685600 369600 687000
rect 371000 685600 372600 687000
rect 374000 685600 375600 687000
rect 377000 685600 378600 687000
rect 380000 685600 381600 687000
rect 383000 685600 384600 687000
rect 386000 685600 387600 687000
rect 389000 685600 390600 687000
rect 392000 685600 393600 687000
rect 395000 685600 396600 687000
rect 398000 685600 399600 687000
rect 401000 685600 402600 687000
rect 404000 685600 405600 687000
rect 407000 685600 408600 687000
rect 410000 685600 411600 687000
rect 413000 685600 414600 687000
rect 416000 685600 417600 687000
rect 419000 685600 420600 687000
rect 422000 685600 423600 687000
rect 425000 685600 426600 687000
rect 428000 685600 429600 687000
rect 431000 685600 432600 687000
rect 434000 685600 435600 687000
rect 437000 685600 438600 687000
rect 440000 685600 441600 687000
rect 443000 685600 444600 687000
rect 446000 685600 447600 687000
rect 449000 685600 450600 687000
rect 452000 685600 453600 687000
rect 455000 685600 456600 687000
rect 458000 685600 459600 687000
rect 461000 685600 462600 687000
rect 464000 685600 465600 687000
rect 467000 685600 468600 687000
rect 470000 685600 471600 687000
rect 473000 685600 474600 687000
rect 476000 685600 477600 687000
rect 479000 685600 480600 687000
rect 482000 685600 483600 687000
rect 485000 685600 486600 687000
rect 488000 685600 489600 687000
rect 491000 685600 492600 687000
rect 494000 685600 495600 687000
rect 497000 685600 498600 687000
rect 500000 685600 501600 687000
rect 503000 685600 504600 687000
rect 506000 685600 507600 687000
rect 509000 685600 510600 687000
rect 512000 685600 513600 687000
rect 515000 685600 516600 687000
rect 518000 685600 519600 687000
rect 521000 685600 522600 687000
rect 524000 685600 525600 687000
rect 5400 682600 7000 684000
rect 9200 682600 10800 684000
rect 14000 682600 15600 684000
rect 17000 682600 18600 684000
rect 20000 682600 21600 684000
rect 23000 682600 24600 684000
rect 26000 682600 27600 684000
rect 29000 682600 30600 684000
rect 32000 682600 33600 684000
rect 35000 682600 36600 684000
rect 38000 682600 39600 684000
rect 41000 682600 42600 684000
rect 44000 682600 45600 684000
rect 47000 682600 48600 684000
rect 50000 682600 51600 684000
rect 53000 682600 54600 684000
rect 56000 682600 57600 684000
rect 59000 682600 60600 684000
rect 62000 682600 63600 684000
rect 65000 682600 66600 684000
rect 68000 682600 69600 684000
rect 71000 682600 72600 684000
rect 74000 682600 75600 684000
rect 77000 682600 78600 684000
rect 80000 682600 81600 684000
rect 83000 682600 84600 684000
rect 86000 682600 87600 684000
rect 89000 682600 90600 684000
rect 92000 682600 93600 684000
rect 95000 682600 96600 684000
rect 98000 682600 99600 684000
rect 101000 682600 102600 684000
rect 104000 682600 105600 684000
rect 107000 682600 108600 684000
rect 110000 682600 111600 684000
rect 113000 682600 114600 684000
rect 116000 682600 117600 684000
rect 119000 682600 120600 684000
rect 122000 682600 123600 684000
rect 125000 682600 126600 684000
rect 128000 682600 129600 684000
rect 131000 682600 132600 684000
rect 134000 682600 135600 684000
rect 137000 682600 138600 684000
rect 140000 682600 141600 684000
rect 143000 682600 144600 684000
rect 146000 682600 147600 684000
rect 149000 682600 150600 684000
rect 152000 682600 153600 684000
rect 155000 682600 156600 684000
rect 158000 682600 159600 684000
rect 161000 682600 162600 684000
rect 164000 682600 165600 684000
rect 167000 682600 168600 684000
rect 170000 682600 171600 684000
rect 173000 682600 174600 684000
rect 176000 682600 177600 684000
rect 179000 682600 180600 684000
rect 182000 682600 183600 684000
rect 185000 682600 186600 684000
rect 188000 682600 189600 684000
rect 191000 682600 192600 684000
rect 194000 682600 195600 684000
rect 197000 682600 198600 684000
rect 200000 682600 201600 684000
rect 203000 682600 204600 684000
rect 206000 682600 207600 684000
rect 209000 682600 210600 684000
rect 212000 682600 213600 684000
rect 215000 682600 216600 684000
rect 218000 682600 219600 684000
rect 221000 682600 222600 684000
rect 224000 682600 225600 684000
rect 227000 682600 228600 684000
rect 230000 682600 231600 684000
rect 233000 682600 234600 684000
rect 236000 682600 237600 684000
rect 239000 682600 240600 684000
rect 242000 682600 243600 684000
rect 245000 682600 246600 684000
rect 248000 682600 249600 684000
rect 251000 682600 252600 684000
rect 254000 682600 255600 684000
rect 257000 682600 258600 684000
rect 260000 682600 261600 684000
rect 263000 682600 264600 684000
rect 266000 682600 267600 684000
rect 269000 682600 270600 684000
rect 272000 682600 273600 684000
rect 275000 682600 276600 684000
rect 278000 682600 279600 684000
rect 281000 682600 282600 684000
rect 284000 682600 285600 684000
rect 287000 682600 288600 684000
rect 290000 682600 291600 684000
rect 293000 682600 294600 684000
rect 296000 682600 297600 684000
rect 299000 682600 300600 684000
rect 302000 682600 303600 684000
rect 305000 682600 306600 684000
rect 308000 682600 309600 684000
rect 311000 682600 312600 684000
rect 314000 682600 315600 684000
rect 317000 682600 318600 684000
rect 320000 682600 321600 684000
rect 323000 682600 324600 684000
rect 326000 682600 327600 684000
rect 329000 682600 330600 684000
rect 332000 682600 333600 684000
rect 335000 682600 336600 684000
rect 338000 682600 339600 684000
rect 341000 682600 342600 684000
rect 344000 682600 345600 684000
rect 347000 682600 348600 684000
rect 350000 682600 351600 684000
rect 353000 682600 354600 684000
rect 356000 682600 357600 684000
rect 359000 682600 360600 684000
rect 362000 682600 363600 684000
rect 365000 682600 366600 684000
rect 368000 682600 369600 684000
rect 371000 682600 372600 684000
rect 374000 682600 375600 684000
rect 377000 682600 378600 684000
rect 380000 682600 381600 684000
rect 383000 682600 384600 684000
rect 386000 682600 387600 684000
rect 389000 682600 390600 684000
rect 392000 682600 393600 684000
rect 395000 682600 396600 684000
rect 398000 682600 399600 684000
rect 401000 682600 402600 684000
rect 404000 682600 405600 684000
rect 407000 682600 408600 684000
rect 410000 682600 411600 684000
rect 413000 682600 414600 684000
rect 416000 682600 417600 684000
rect 419000 682600 420600 684000
rect 422000 682600 423600 684000
rect 425000 682600 426600 684000
rect 428000 682600 429600 684000
rect 431000 682600 432600 684000
rect 434000 682600 435600 684000
rect 437000 682600 438600 684000
rect 440000 682600 441600 684000
rect 443000 682600 444600 684000
rect 446000 682600 447600 684000
rect 449000 682600 450600 684000
rect 452000 682600 453600 684000
rect 455000 682600 456600 684000
rect 458000 682600 459600 684000
rect 461000 682600 462600 684000
rect 464000 682600 465600 684000
rect 467000 682600 468600 684000
rect 470000 682600 471600 684000
rect 473000 682600 474600 684000
rect 476000 682600 477600 684000
rect 479000 682600 480600 684000
rect 482000 682600 483600 684000
rect 485000 682600 486600 684000
rect 488000 682600 489600 684000
rect 491000 682600 492600 684000
rect 494000 682600 495600 684000
rect 497000 682600 498600 684000
rect 500000 682600 501600 684000
rect 503000 682600 504600 684000
rect 506000 682600 507600 684000
rect 509000 682600 510600 684000
rect 512000 682600 513600 684000
rect 515000 682600 516600 684000
rect 518000 682600 519600 684000
rect 521000 682600 522600 684000
rect 524000 682600 525600 684000
rect 5400 679600 7000 681000
rect 9200 679600 10800 681000
rect 14000 679600 15600 681000
rect 5400 676600 7000 678000
rect 9200 676600 10800 678000
rect 14000 676600 15600 678000
rect 580470 678030 581910 682990
rect 5400 673600 7000 675000
rect 9200 673600 10800 675000
rect 14000 673600 15600 675000
rect 5400 670600 7000 672000
rect 9200 670600 10800 672000
rect 14000 670600 15600 672000
rect 5400 667600 7000 669000
rect 9200 667600 10800 669000
rect 14000 667600 15600 669000
rect 512660 667690 513650 668160
rect 5400 664600 7000 666000
rect 9200 664600 10800 666000
rect 14000 664600 15600 666000
rect 512420 664910 514020 665220
rect 520580 664340 526480 669740
rect 5400 661600 7000 663000
rect 9200 661600 10800 663000
rect 14000 661600 15600 663000
rect 5400 658600 7000 660000
rect 9200 658600 10800 660000
rect 14000 658600 15600 660000
rect 5400 655600 7000 657000
rect 9200 655600 10800 657000
rect 14000 655600 15600 657000
rect 5400 652600 7000 654000
rect 9200 652600 10800 654000
rect 14000 652600 15600 654000
rect 503480 652270 503670 653460
rect 5400 649600 7000 651000
rect 9200 649600 10800 651000
rect 14000 649600 15600 651000
rect 5400 646600 7000 648000
rect 9200 646600 10800 648000
rect 14000 646600 15600 648000
rect 5400 643600 7000 645000
rect 9200 643600 10800 645000
rect 14000 643600 15600 645000
rect 5400 640600 7000 642000
rect 9200 640600 10800 642000
rect 14000 640600 15600 642000
rect 5400 637600 7000 639000
rect 9200 637600 10800 639000
rect 14000 637600 15600 639000
rect 5400 634600 7000 636000
rect 9200 634600 10800 636000
rect 14000 634600 15600 636000
rect 5400 631600 7000 633000
rect 9200 631600 10800 633000
rect 14000 631600 15600 633000
rect 5400 628600 7000 630000
rect 9200 628600 10800 630000
rect 14000 628600 15600 630000
rect 5400 625600 7000 627000
rect 9200 625600 10800 627000
rect 14000 625600 15600 627000
rect 5400 622600 7000 624000
rect 9200 622600 10800 624000
rect 14000 622600 15600 624000
rect 5400 619600 7000 621000
rect 9200 619600 10800 621000
rect 14000 619600 15600 621000
rect 5400 616600 7000 618000
rect 9200 616600 10800 618000
rect 14000 616600 15600 618000
rect 520780 641340 526680 646740
rect 576690 630020 583530 644270
rect 520580 617740 526580 623040
rect 5400 613600 7000 615000
rect 9200 613600 10800 615000
rect 14000 613600 15600 615000
rect 5400 610600 7000 612000
rect 9200 610600 10800 612000
rect 14000 610600 15600 612000
rect 5400 607600 7000 609000
rect 9200 607600 10800 609000
rect 14000 607600 15600 609000
rect 5400 604600 7000 606000
rect 9200 604600 10800 606000
rect 14000 604600 15600 606000
rect 5400 601600 7000 603000
rect 9200 601600 10800 603000
rect 14000 601600 15600 603000
rect 5400 598600 7000 600000
rect 9200 598600 10800 600000
rect 14000 598600 15600 600000
rect 5400 595600 7000 597000
rect 9200 595600 10800 597000
rect 14000 595600 15600 597000
rect 5400 592600 7000 594000
rect 9200 592600 10800 594000
rect 14000 592600 15600 594000
rect 5400 589600 7000 591000
rect 9200 589600 10800 591000
rect 14000 589600 15600 591000
rect 5400 586600 7000 588000
rect 9200 586600 10800 588000
rect 14000 586600 15600 588000
rect 5400 583600 7000 585000
rect 9200 583600 10800 585000
rect 14000 583600 15600 585000
rect 5400 580600 7000 582000
rect 9200 580600 10800 582000
rect 14000 580600 15600 582000
rect 577730 580390 583180 583570
rect 5400 577600 7000 579000
rect 9200 577600 10800 579000
rect 14000 577600 15600 579000
rect 5400 574600 7000 576000
rect 9200 574600 10800 576000
rect 14000 574600 15600 576000
rect 5400 571600 7000 573000
rect 9200 571600 10800 573000
rect 14000 571600 15600 573000
rect 504870 572030 505860 572500
rect 5400 568600 7000 570000
rect 9200 568600 10800 570000
rect 14000 568600 15600 570000
rect 504630 569250 506230 569560
rect 512590 568680 518490 574080
rect 557460 572160 558450 572630
rect 557220 569380 558820 569690
rect 565180 568810 571080 574210
rect 5400 565600 7000 567000
rect 9200 565600 10800 567000
rect 14000 565600 15600 567000
rect 870 549250 2600 564320
rect 4400 563000 6000 564400
rect 7200 563000 8800 564400
rect 9800 563000 11400 564400
rect 12800 563000 14400 564400
rect 15600 563000 17200 564400
rect 4400 560000 6000 561400
rect 7200 560000 8800 561400
rect 9800 560000 11400 561400
rect 12800 560000 14400 561400
rect 15600 560000 17200 561400
rect 4400 556800 6000 558200
rect 7200 556800 8800 558200
rect 9800 556800 11400 558200
rect 12800 556800 14400 558200
rect 15600 556800 17200 558200
rect 495490 556610 495680 557800
rect 4400 554400 6000 555800
rect 7200 554400 8800 555800
rect 9800 554400 11400 555800
rect 12800 554400 14400 555800
rect 15600 554400 17200 555800
rect 4400 551800 6000 553200
rect 7200 551800 8800 553200
rect 9800 551800 11400 553200
rect 12800 551800 14400 553200
rect 15600 551800 17200 553200
rect 16000 551600 16600 551800
rect 4400 549200 6000 550600
rect 7200 549200 8800 550600
rect 9800 549200 11400 550600
rect 12800 549200 14400 550600
rect 15600 549200 17200 550600
rect 16000 548600 16600 549200
rect 6920 534720 7200 536700
rect 8420 534720 8700 536700
rect 548080 556740 548270 557930
rect 512790 545680 518690 551080
rect 565380 545810 571280 551210
rect 512590 522080 518590 527380
rect 565180 522210 571180 527510
rect 300 511100 2350 512460
rect 553320 496420 554510 496610
rect 565960 485870 566270 487470
rect 580590 493390 582340 495690
rect 568740 486240 569210 487230
rect 518790 473510 524090 479510
rect 542390 473410 547790 479310
rect 565390 473610 570790 479510
rect 330 467850 2380 469210
rect 576750 448670 578500 450970
rect 400 423400 1800 424600
rect 571720 405820 577750 407140
rect 400 380100 1800 381300
rect 574000 363400 574600 364800
rect 575800 363400 576000 365000
rect 576800 363400 577400 364800
rect 578600 363400 578800 365000
rect 572600 361200 573400 361400
rect 573800 361200 574600 361400
rect 572600 360800 573400 361000
rect 573800 360800 574600 361000
rect 572600 360400 573400 360600
rect 573800 360400 574600 360600
rect 572600 360000 573400 360200
rect 573800 360000 574600 360200
rect 572600 359600 573400 359800
rect 573800 359600 574600 359800
rect 572600 359200 573400 359400
rect 573800 359200 574600 359400
rect 579150 359440 582190 360800
rect 572600 358800 573400 359000
rect 573800 358800 574600 359000
rect 572600 358400 573400 358600
rect 573800 358400 574600 358600
rect 572600 358000 573400 358200
rect 573800 358000 574600 358200
rect 572600 357600 573400 357800
rect 573800 357600 574600 357800
rect 572600 357200 573400 357400
rect 573800 357200 574600 357400
rect 572600 356800 573400 357000
rect 573800 356800 574600 357000
rect 572600 356400 573400 356600
rect 573800 356400 574600 356600
rect 572600 356000 573400 356200
rect 573800 356000 574600 356200
rect 572600 355600 573400 355800
rect 573800 355600 574600 355800
rect 572600 355200 573400 355400
rect 573800 355200 574600 355400
rect 572600 354800 573400 355000
rect 573800 354800 574600 355000
rect 572600 354400 573400 354600
rect 573800 354400 574600 354600
rect 572600 354000 573400 354200
rect 573800 354000 574600 354200
rect 6123 343490 6313 344680
rect 400 336900 1800 338100
rect 2930 324813 3240 326413
rect 5710 325183 6180 326173
rect 400 294900 1800 296100
rect 400 251800 1800 253000
rect 700 163110 2330 177370
rect 576980 314100 579620 315490
rect 573690 269790 579290 270990
rect 572040 216420 572230 217610
rect 579460 198160 580960 201000
rect 579500 189900 580900 198160
rect 576400 167200 579400 175500
rect 573200 151830 576200 152000
rect 573150 148990 576200 151830
rect 573200 143700 576200 148990
rect 570880 130770 577350 130820
rect 400 124300 1800 125500
rect 570850 123400 577320 130770
rect 577320 123400 577350 130770
<< metal3 >>
rect 16194 703660 21194 704800
rect 15390 703180 21970 703660
rect 68194 703470 73194 704800
rect 15390 701230 15690 703180
rect 21540 701230 21970 703180
rect 67560 703110 73630 703470
rect 67560 701700 67850 703110
rect 73380 701700 73630 703110
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702990 232594 704800
rect 227594 702520 233090 702990
rect 227594 702300 228670 702520
rect 222800 702000 224600 702300
rect 67560 701540 73630 701700
rect 15390 700950 21970 701230
rect 214000 700200 224600 702000
rect 214000 693800 219400 700200
rect 222800 700000 224600 700200
rect 225200 699600 227200 702300
rect 228240 701850 228670 702300
rect 232530 701850 233090 702520
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702880 334294 704800
rect 329294 702410 334900 702880
rect 329294 702300 330480 702410
rect 324400 702000 326200 702300
rect 228240 701380 233090 701850
rect 222200 698800 227200 699600
rect 222200 698000 222600 698800
rect 226600 698000 227200 698800
rect 222200 697600 227200 698000
rect 222200 696800 222600 697600
rect 226600 696800 227200 697600
rect 222200 696400 227200 696800
rect 222200 695600 222600 696400
rect 226600 695600 227200 696400
rect 222200 695400 227200 695600
rect 316200 700000 326200 702000
rect 316200 693800 322200 700000
rect 326800 699600 328800 702300
rect 330050 701740 330480 702300
rect 334340 701740 334900 702410
rect 413394 702300 418394 704800
rect 465394 703610 470394 704800
rect 510594 703780 515394 704800
rect 520594 703780 525394 704800
rect 330050 701270 334900 701740
rect 463110 701590 471840 703610
rect 510594 703440 525450 703780
rect 510594 702340 510880 703440
rect 323800 698800 328800 699600
rect 463110 699400 463720 701590
rect 471140 699400 471840 701590
rect 510600 700600 510880 702340
rect 463110 698980 471840 699400
rect 323800 698000 324200 698800
rect 328200 698000 328800 698800
rect 323800 697600 328800 698000
rect 323800 696800 324200 697600
rect 328200 696800 328800 697600
rect 323800 696400 328800 696800
rect 323800 695600 324200 696400
rect 328200 695600 328800 696400
rect 323800 695400 328800 695600
rect 510000 696600 510880 700600
rect 525130 700600 525450 703440
rect 566594 702930 571594 704800
rect 565960 701120 573480 702930
rect 525130 696600 526600 700600
rect 565960 699450 566440 701120
rect 573030 699450 573480 701120
rect 565960 698710 573480 699450
rect 510000 693800 526600 696600
rect 4400 693000 526600 693800
rect 4400 691600 5400 693000
rect 7000 691600 9200 693000
rect 10800 691600 14000 693000
rect 15600 691600 17000 693000
rect 18600 691600 20000 693000
rect 21600 691600 23000 693000
rect 24600 691600 26000 693000
rect 27600 691600 29000 693000
rect 30600 691600 32000 693000
rect 33600 691600 35000 693000
rect 36600 691600 38000 693000
rect 39600 691600 41000 693000
rect 42600 691600 44000 693000
rect 45600 691600 47000 693000
rect 48600 691600 50000 693000
rect 51600 691600 53000 693000
rect 54600 691600 56000 693000
rect 57600 691600 59000 693000
rect 60600 691600 62000 693000
rect 63600 691600 65000 693000
rect 66600 691600 68000 693000
rect 69600 691600 71000 693000
rect 72600 691600 74000 693000
rect 75600 691600 77000 693000
rect 78600 691600 80000 693000
rect 81600 691600 83000 693000
rect 84600 691600 86000 693000
rect 87600 691600 89000 693000
rect 90600 691600 92000 693000
rect 93600 691600 95000 693000
rect 96600 691600 98000 693000
rect 99600 691600 101000 693000
rect 102600 691600 104000 693000
rect 105600 691600 107000 693000
rect 108600 691600 110000 693000
rect 111600 691600 113000 693000
rect 114600 691600 116000 693000
rect 117600 691600 119000 693000
rect 120600 691600 122000 693000
rect 123600 691600 125000 693000
rect 126600 691600 128000 693000
rect 129600 691600 131000 693000
rect 132600 691600 134000 693000
rect 135600 691600 137000 693000
rect 138600 691600 140000 693000
rect 141600 691600 143000 693000
rect 144600 691600 146000 693000
rect 147600 691600 149000 693000
rect 150600 691600 152000 693000
rect 153600 691600 155000 693000
rect 156600 691600 158000 693000
rect 159600 691600 161000 693000
rect 162600 691600 164000 693000
rect 165600 691600 167000 693000
rect 168600 691600 170000 693000
rect 171600 691600 173000 693000
rect 174600 691600 176000 693000
rect 177600 691600 179000 693000
rect 180600 691600 182000 693000
rect 183600 691600 185000 693000
rect 186600 691600 188000 693000
rect 189600 691600 191000 693000
rect 192600 691600 194000 693000
rect 195600 691600 197000 693000
rect 198600 691600 200000 693000
rect 201600 691600 203000 693000
rect 204600 691600 206000 693000
rect 207600 691600 209000 693000
rect 210600 691600 212000 693000
rect 213600 691600 215000 693000
rect 216600 691600 218000 693000
rect 219600 691600 221000 693000
rect 222600 691600 224000 693000
rect 225600 691600 227000 693000
rect 228600 691600 230000 693000
rect 231600 691600 233000 693000
rect 234600 691600 236000 693000
rect 237600 691600 239000 693000
rect 240600 691600 242000 693000
rect 243600 691600 245000 693000
rect 246600 691600 248000 693000
rect 249600 691600 251000 693000
rect 252600 691600 254000 693000
rect 255600 691600 257000 693000
rect 258600 691600 260000 693000
rect 261600 691600 263000 693000
rect 264600 691600 266000 693000
rect 267600 691600 269000 693000
rect 270600 691600 272000 693000
rect 273600 691600 275000 693000
rect 276600 691600 278000 693000
rect 279600 691600 281000 693000
rect 282600 691600 284000 693000
rect 285600 691600 287000 693000
rect 288600 691600 290000 693000
rect 291600 691600 293000 693000
rect 294600 691600 296000 693000
rect 297600 691600 299000 693000
rect 300600 691600 302000 693000
rect 303600 691600 305000 693000
rect 306600 691600 308000 693000
rect 309600 691600 311000 693000
rect 312600 691600 314000 693000
rect 315600 691600 317000 693000
rect 318600 691600 320000 693000
rect 321600 691600 323000 693000
rect 324600 691600 326000 693000
rect 327600 691600 329000 693000
rect 330600 691600 332000 693000
rect 333600 691600 335000 693000
rect 336600 691600 338000 693000
rect 339600 691600 341000 693000
rect 342600 691600 344000 693000
rect 345600 691600 347000 693000
rect 348600 691600 350000 693000
rect 351600 691600 353000 693000
rect 354600 691600 356000 693000
rect 357600 691600 359000 693000
rect 360600 691600 362000 693000
rect 363600 691600 365000 693000
rect 366600 691600 368000 693000
rect 369600 691600 371000 693000
rect 372600 691600 374000 693000
rect 375600 691600 377000 693000
rect 378600 691600 380000 693000
rect 381600 691600 383000 693000
rect 384600 691600 386000 693000
rect 387600 691600 389000 693000
rect 390600 691600 392000 693000
rect 393600 691600 395000 693000
rect 396600 691600 398000 693000
rect 399600 691600 401000 693000
rect 402600 691600 404000 693000
rect 405600 691600 407000 693000
rect 408600 691600 410000 693000
rect 411600 691600 413000 693000
rect 414600 691600 416000 693000
rect 417600 691600 419000 693000
rect 420600 691600 422000 693000
rect 423600 691600 425000 693000
rect 426600 691600 428000 693000
rect 429600 691600 431000 693000
rect 432600 691600 434000 693000
rect 435600 691600 437000 693000
rect 438600 691600 440000 693000
rect 441600 691600 443000 693000
rect 444600 691600 446000 693000
rect 447600 691600 449000 693000
rect 450600 691600 452000 693000
rect 453600 691600 455000 693000
rect 456600 691600 458000 693000
rect 459600 691600 461000 693000
rect 462600 691600 464000 693000
rect 465600 691600 467000 693000
rect 468600 691600 470000 693000
rect 471600 691600 473000 693000
rect 474600 691600 476000 693000
rect 477600 691600 479000 693000
rect 480600 691600 482000 693000
rect 483600 691600 485000 693000
rect 486600 691600 488000 693000
rect 489600 691600 491000 693000
rect 492600 691600 494000 693000
rect 495600 691600 497000 693000
rect 498600 691600 500000 693000
rect 501600 691600 503000 693000
rect 504600 691600 506000 693000
rect 507600 691600 509000 693000
rect 510600 691600 512000 693000
rect 513600 691600 515000 693000
rect 516600 691600 518000 693000
rect 519600 691600 521000 693000
rect 522600 691600 524000 693000
rect 525600 691600 526600 693000
rect 4400 690000 526600 691600
rect 4400 688600 5400 690000
rect 7000 688600 9200 690000
rect 10800 688600 14000 690000
rect 15600 688600 17000 690000
rect 18600 688600 20000 690000
rect 21600 688600 23000 690000
rect 24600 688600 26000 690000
rect 27600 688600 29000 690000
rect 30600 688600 32000 690000
rect 33600 688600 35000 690000
rect 36600 688600 38000 690000
rect 39600 688600 41000 690000
rect 42600 688600 44000 690000
rect 45600 688600 47000 690000
rect 48600 688600 50000 690000
rect 51600 688600 53000 690000
rect 54600 688600 56000 690000
rect 57600 688600 59000 690000
rect 60600 688600 62000 690000
rect 63600 688600 65000 690000
rect 66600 688600 68000 690000
rect 69600 688600 71000 690000
rect 72600 688600 74000 690000
rect 75600 688600 77000 690000
rect 78600 688600 80000 690000
rect 81600 688600 83000 690000
rect 84600 688600 86000 690000
rect 87600 688600 89000 690000
rect 90600 688600 92000 690000
rect 93600 688600 95000 690000
rect 96600 688600 98000 690000
rect 99600 688600 101000 690000
rect 102600 688600 104000 690000
rect 105600 688600 107000 690000
rect 108600 688600 110000 690000
rect 111600 688600 113000 690000
rect 114600 688600 116000 690000
rect 117600 688600 119000 690000
rect 120600 688600 122000 690000
rect 123600 688600 125000 690000
rect 126600 688600 128000 690000
rect 129600 688600 131000 690000
rect 132600 688600 134000 690000
rect 135600 688600 137000 690000
rect 138600 688600 140000 690000
rect 141600 688600 143000 690000
rect 144600 688600 146000 690000
rect 147600 688600 149000 690000
rect 150600 688600 152000 690000
rect 153600 688600 155000 690000
rect 156600 688600 158000 690000
rect 159600 688600 161000 690000
rect 162600 688600 164000 690000
rect 165600 688600 167000 690000
rect 168600 688600 170000 690000
rect 171600 688600 173000 690000
rect 174600 688600 176000 690000
rect 177600 688600 179000 690000
rect 180600 688600 182000 690000
rect 183600 688600 185000 690000
rect 186600 688600 188000 690000
rect 189600 688600 191000 690000
rect 192600 688600 194000 690000
rect 195600 688600 197000 690000
rect 198600 688600 200000 690000
rect 201600 688600 203000 690000
rect 204600 688600 206000 690000
rect 207600 688600 209000 690000
rect 210600 688600 212000 690000
rect 213600 688600 215000 690000
rect 216600 688600 218000 690000
rect 219600 688600 221000 690000
rect 222600 688600 224000 690000
rect 225600 688600 227000 690000
rect 228600 688600 230000 690000
rect 231600 688600 233000 690000
rect 234600 688600 236000 690000
rect 237600 688600 239000 690000
rect 240600 688600 242000 690000
rect 243600 688600 245000 690000
rect 246600 688600 248000 690000
rect 249600 688600 251000 690000
rect 252600 688600 254000 690000
rect 255600 688600 257000 690000
rect 258600 688600 260000 690000
rect 261600 688600 263000 690000
rect 264600 688600 266000 690000
rect 267600 688600 269000 690000
rect 270600 688600 272000 690000
rect 273600 688600 275000 690000
rect 276600 688600 278000 690000
rect 279600 688600 281000 690000
rect 282600 688600 284000 690000
rect 285600 688600 287000 690000
rect 288600 688600 290000 690000
rect 291600 688600 293000 690000
rect 294600 688600 296000 690000
rect 297600 688600 299000 690000
rect 300600 688600 302000 690000
rect 303600 688600 305000 690000
rect 306600 688600 308000 690000
rect 309600 688600 311000 690000
rect 312600 688600 314000 690000
rect 315600 688600 317000 690000
rect 318600 688600 320000 690000
rect 321600 688600 323000 690000
rect 324600 688600 326000 690000
rect 327600 688600 329000 690000
rect 330600 688600 332000 690000
rect 333600 688600 335000 690000
rect 336600 688600 338000 690000
rect 339600 688600 341000 690000
rect 342600 688600 344000 690000
rect 345600 688600 347000 690000
rect 348600 688600 350000 690000
rect 351600 688600 353000 690000
rect 354600 688600 356000 690000
rect 357600 688600 359000 690000
rect 360600 688600 362000 690000
rect 363600 688600 365000 690000
rect 366600 688600 368000 690000
rect 369600 688600 371000 690000
rect 372600 688600 374000 690000
rect 375600 688600 377000 690000
rect 378600 688600 380000 690000
rect 381600 688600 383000 690000
rect 384600 688600 386000 690000
rect 387600 688600 389000 690000
rect 390600 688600 392000 690000
rect 393600 688600 395000 690000
rect 396600 688600 398000 690000
rect 399600 688600 401000 690000
rect 402600 688600 404000 690000
rect 405600 688600 407000 690000
rect 408600 688600 410000 690000
rect 411600 688600 413000 690000
rect 414600 688600 416000 690000
rect 417600 688600 419000 690000
rect 420600 688600 422000 690000
rect 423600 688600 425000 690000
rect 426600 688600 428000 690000
rect 429600 688600 431000 690000
rect 432600 688600 434000 690000
rect 435600 688600 437000 690000
rect 438600 688600 440000 690000
rect 441600 688600 443000 690000
rect 444600 688600 446000 690000
rect 447600 688600 449000 690000
rect 450600 688600 452000 690000
rect 453600 688600 455000 690000
rect 456600 688600 458000 690000
rect 459600 688600 461000 690000
rect 462600 688600 464000 690000
rect 465600 688600 467000 690000
rect 468600 688600 470000 690000
rect 471600 688600 473000 690000
rect 474600 688600 476000 690000
rect 477600 688600 479000 690000
rect 480600 688600 482000 690000
rect 483600 688600 485000 690000
rect 486600 688600 488000 690000
rect 489600 688600 491000 690000
rect 492600 688600 494000 690000
rect 495600 688600 497000 690000
rect 498600 688600 500000 690000
rect 501600 688600 503000 690000
rect 504600 688600 506000 690000
rect 507600 688600 509000 690000
rect 510600 688600 512000 690000
rect 513600 688600 515000 690000
rect 516600 688600 518000 690000
rect 519600 688600 521000 690000
rect 522600 688600 524000 690000
rect 525600 688600 526600 690000
rect 4400 687000 526600 688600
rect 930 685550 3360 685890
rect 930 685242 1340 685550
rect -800 680242 1340 685242
rect 930 679860 1340 680242
rect 3090 679860 3360 685550
rect 930 679660 3360 679860
rect 4400 685600 5400 687000
rect 7000 685600 9200 687000
rect 10800 685600 14000 687000
rect 15600 685600 17000 687000
rect 18600 685600 20000 687000
rect 21600 685600 23000 687000
rect 24600 685600 26000 687000
rect 27600 685600 29000 687000
rect 30600 685600 32000 687000
rect 33600 685600 35000 687000
rect 36600 685600 38000 687000
rect 39600 685600 41000 687000
rect 42600 685600 44000 687000
rect 45600 685600 47000 687000
rect 48600 685600 50000 687000
rect 51600 685600 53000 687000
rect 54600 685600 56000 687000
rect 57600 685600 59000 687000
rect 60600 685600 62000 687000
rect 63600 685600 65000 687000
rect 66600 685600 68000 687000
rect 69600 685600 71000 687000
rect 72600 685600 74000 687000
rect 75600 685600 77000 687000
rect 78600 685600 80000 687000
rect 81600 685600 83000 687000
rect 84600 685600 86000 687000
rect 87600 685600 89000 687000
rect 90600 685600 92000 687000
rect 93600 685600 95000 687000
rect 96600 685600 98000 687000
rect 99600 685600 101000 687000
rect 102600 685600 104000 687000
rect 105600 685600 107000 687000
rect 108600 685600 110000 687000
rect 111600 685600 113000 687000
rect 114600 685600 116000 687000
rect 117600 685600 119000 687000
rect 120600 685600 122000 687000
rect 123600 685600 125000 687000
rect 126600 685600 128000 687000
rect 129600 685600 131000 687000
rect 132600 685600 134000 687000
rect 135600 685600 137000 687000
rect 138600 685600 140000 687000
rect 141600 685600 143000 687000
rect 144600 685600 146000 687000
rect 147600 685600 149000 687000
rect 150600 685600 152000 687000
rect 153600 685600 155000 687000
rect 156600 685600 158000 687000
rect 159600 685600 161000 687000
rect 162600 685600 164000 687000
rect 165600 685600 167000 687000
rect 168600 685600 170000 687000
rect 171600 685600 173000 687000
rect 174600 685600 176000 687000
rect 177600 685600 179000 687000
rect 180600 685600 182000 687000
rect 183600 685600 185000 687000
rect 186600 685600 188000 687000
rect 189600 685600 191000 687000
rect 192600 685600 194000 687000
rect 195600 685600 197000 687000
rect 198600 685600 200000 687000
rect 201600 685600 203000 687000
rect 204600 685600 206000 687000
rect 207600 685600 209000 687000
rect 210600 685600 212000 687000
rect 213600 685600 215000 687000
rect 216600 685600 218000 687000
rect 219600 685600 221000 687000
rect 222600 685600 224000 687000
rect 225600 685600 227000 687000
rect 228600 685600 230000 687000
rect 231600 685600 233000 687000
rect 234600 685600 236000 687000
rect 237600 685600 239000 687000
rect 240600 685600 242000 687000
rect 243600 685600 245000 687000
rect 246600 685600 248000 687000
rect 249600 685600 251000 687000
rect 252600 685600 254000 687000
rect 255600 685600 257000 687000
rect 258600 685600 260000 687000
rect 261600 685600 263000 687000
rect 264600 685600 266000 687000
rect 267600 685600 269000 687000
rect 270600 685600 272000 687000
rect 273600 685600 275000 687000
rect 276600 685600 278000 687000
rect 279600 685600 281000 687000
rect 282600 685600 284000 687000
rect 285600 685600 287000 687000
rect 288600 685600 290000 687000
rect 291600 685600 293000 687000
rect 294600 685600 296000 687000
rect 297600 685600 299000 687000
rect 300600 685600 302000 687000
rect 303600 685600 305000 687000
rect 306600 685600 308000 687000
rect 309600 685600 311000 687000
rect 312600 685600 314000 687000
rect 315600 685600 317000 687000
rect 318600 685600 320000 687000
rect 321600 685600 323000 687000
rect 324600 685600 326000 687000
rect 327600 685600 329000 687000
rect 330600 685600 332000 687000
rect 333600 685600 335000 687000
rect 336600 685600 338000 687000
rect 339600 685600 341000 687000
rect 342600 685600 344000 687000
rect 345600 685600 347000 687000
rect 348600 685600 350000 687000
rect 351600 685600 353000 687000
rect 354600 685600 356000 687000
rect 357600 685600 359000 687000
rect 360600 685600 362000 687000
rect 363600 685600 365000 687000
rect 366600 685600 368000 687000
rect 369600 685600 371000 687000
rect 372600 685600 374000 687000
rect 375600 685600 377000 687000
rect 378600 685600 380000 687000
rect 381600 685600 383000 687000
rect 384600 685600 386000 687000
rect 387600 685600 389000 687000
rect 390600 685600 392000 687000
rect 393600 685600 395000 687000
rect 396600 685600 398000 687000
rect 399600 685600 401000 687000
rect 402600 685600 404000 687000
rect 405600 685600 407000 687000
rect 408600 685600 410000 687000
rect 411600 685600 413000 687000
rect 414600 685600 416000 687000
rect 417600 685600 419000 687000
rect 420600 685600 422000 687000
rect 423600 685600 425000 687000
rect 426600 685600 428000 687000
rect 429600 685600 431000 687000
rect 432600 685600 434000 687000
rect 435600 685600 437000 687000
rect 438600 685600 440000 687000
rect 441600 685600 443000 687000
rect 444600 685600 446000 687000
rect 447600 685600 449000 687000
rect 450600 685600 452000 687000
rect 453600 685600 455000 687000
rect 456600 685600 458000 687000
rect 459600 685600 461000 687000
rect 462600 685600 464000 687000
rect 465600 685600 467000 687000
rect 468600 685600 470000 687000
rect 471600 685600 473000 687000
rect 474600 685600 476000 687000
rect 477600 685600 479000 687000
rect 480600 685600 482000 687000
rect 483600 685600 485000 687000
rect 486600 685600 488000 687000
rect 489600 685600 491000 687000
rect 492600 685600 494000 687000
rect 495600 685600 497000 687000
rect 498600 685600 500000 687000
rect 501600 685600 503000 687000
rect 504600 685600 506000 687000
rect 507600 685600 509000 687000
rect 510600 685600 512000 687000
rect 513600 685600 515000 687000
rect 516600 685600 518000 687000
rect 519600 685600 521000 687000
rect 522600 685600 524000 687000
rect 525600 685600 526600 687000
rect 4400 684000 526600 685600
rect 4400 682600 5400 684000
rect 7000 682600 9200 684000
rect 10800 682600 14000 684000
rect 15600 682600 17000 684000
rect 18600 682600 20000 684000
rect 21600 682600 23000 684000
rect 24600 682600 26000 684000
rect 27600 682600 29000 684000
rect 30600 682600 32000 684000
rect 33600 682600 35000 684000
rect 36600 682600 38000 684000
rect 39600 682600 41000 684000
rect 42600 682600 44000 684000
rect 45600 682600 47000 684000
rect 48600 682600 50000 684000
rect 51600 682600 53000 684000
rect 54600 682600 56000 684000
rect 57600 682600 59000 684000
rect 60600 682600 62000 684000
rect 63600 682600 65000 684000
rect 66600 682600 68000 684000
rect 69600 682600 71000 684000
rect 72600 682600 74000 684000
rect 75600 682600 77000 684000
rect 78600 682600 80000 684000
rect 81600 682600 83000 684000
rect 84600 682600 86000 684000
rect 87600 682600 89000 684000
rect 90600 682600 92000 684000
rect 93600 682600 95000 684000
rect 96600 682600 98000 684000
rect 99600 682600 101000 684000
rect 102600 682600 104000 684000
rect 105600 682600 107000 684000
rect 108600 682600 110000 684000
rect 111600 682600 113000 684000
rect 114600 682600 116000 684000
rect 117600 682600 119000 684000
rect 120600 682600 122000 684000
rect 123600 682600 125000 684000
rect 126600 682600 128000 684000
rect 129600 682600 131000 684000
rect 132600 682600 134000 684000
rect 135600 682600 137000 684000
rect 138600 682600 140000 684000
rect 141600 682600 143000 684000
rect 144600 682600 146000 684000
rect 147600 682600 149000 684000
rect 150600 682600 152000 684000
rect 153600 682600 155000 684000
rect 156600 682600 158000 684000
rect 159600 682600 161000 684000
rect 162600 682600 164000 684000
rect 165600 682600 167000 684000
rect 168600 682600 170000 684000
rect 171600 682600 173000 684000
rect 174600 682600 176000 684000
rect 177600 682600 179000 684000
rect 180600 682600 182000 684000
rect 183600 682600 185000 684000
rect 186600 682600 188000 684000
rect 189600 682600 191000 684000
rect 192600 682600 194000 684000
rect 195600 682600 197000 684000
rect 198600 682600 200000 684000
rect 201600 682600 203000 684000
rect 204600 682600 206000 684000
rect 207600 682600 209000 684000
rect 210600 682600 212000 684000
rect 213600 682600 215000 684000
rect 216600 682600 218000 684000
rect 219600 682600 221000 684000
rect 222600 682600 224000 684000
rect 225600 682600 227000 684000
rect 228600 682600 230000 684000
rect 231600 682600 233000 684000
rect 234600 682600 236000 684000
rect 237600 682600 239000 684000
rect 240600 682600 242000 684000
rect 243600 682600 245000 684000
rect 246600 682600 248000 684000
rect 249600 682600 251000 684000
rect 252600 682600 254000 684000
rect 255600 682600 257000 684000
rect 258600 682600 260000 684000
rect 261600 682600 263000 684000
rect 264600 682600 266000 684000
rect 267600 682600 269000 684000
rect 270600 682600 272000 684000
rect 273600 682600 275000 684000
rect 276600 682600 278000 684000
rect 279600 682600 281000 684000
rect 282600 682600 284000 684000
rect 285600 682600 287000 684000
rect 288600 682600 290000 684000
rect 291600 682600 293000 684000
rect 294600 682600 296000 684000
rect 297600 682600 299000 684000
rect 300600 682600 302000 684000
rect 303600 682600 305000 684000
rect 306600 682600 308000 684000
rect 309600 682600 311000 684000
rect 312600 682600 314000 684000
rect 315600 682600 317000 684000
rect 318600 682600 320000 684000
rect 321600 682600 323000 684000
rect 324600 682600 326000 684000
rect 327600 682600 329000 684000
rect 330600 682600 332000 684000
rect 333600 682600 335000 684000
rect 336600 682600 338000 684000
rect 339600 682600 341000 684000
rect 342600 682600 344000 684000
rect 345600 682600 347000 684000
rect 348600 682600 350000 684000
rect 351600 682600 353000 684000
rect 354600 682600 356000 684000
rect 357600 682600 359000 684000
rect 360600 682600 362000 684000
rect 363600 682600 365000 684000
rect 366600 682600 368000 684000
rect 369600 682600 371000 684000
rect 372600 682600 374000 684000
rect 375600 682600 377000 684000
rect 378600 682600 380000 684000
rect 381600 682600 383000 684000
rect 384600 682600 386000 684000
rect 387600 682600 389000 684000
rect 390600 682600 392000 684000
rect 393600 682600 395000 684000
rect 396600 682600 398000 684000
rect 399600 682600 401000 684000
rect 402600 682600 404000 684000
rect 405600 682600 407000 684000
rect 408600 682600 410000 684000
rect 411600 682600 413000 684000
rect 414600 682600 416000 684000
rect 417600 682600 419000 684000
rect 420600 682600 422000 684000
rect 423600 682600 425000 684000
rect 426600 682600 428000 684000
rect 429600 682600 431000 684000
rect 432600 682600 434000 684000
rect 435600 682600 437000 684000
rect 438600 682600 440000 684000
rect 441600 682600 443000 684000
rect 444600 682600 446000 684000
rect 447600 682600 449000 684000
rect 450600 682600 452000 684000
rect 453600 682600 455000 684000
rect 456600 682600 458000 684000
rect 459600 682600 461000 684000
rect 462600 682600 464000 684000
rect 465600 682600 467000 684000
rect 468600 682600 470000 684000
rect 471600 682600 473000 684000
rect 474600 682600 476000 684000
rect 477600 682600 479000 684000
rect 480600 682600 482000 684000
rect 483600 682600 485000 684000
rect 486600 682600 488000 684000
rect 489600 682600 491000 684000
rect 492600 682600 494000 684000
rect 495600 682600 497000 684000
rect 498600 682600 500000 684000
rect 501600 682600 503000 684000
rect 504600 682600 506000 684000
rect 507600 682600 509000 684000
rect 510600 682600 512000 684000
rect 513600 682600 515000 684000
rect 516600 682600 518000 684000
rect 519600 682600 521000 684000
rect 522600 682600 524000 684000
rect 525600 682600 526600 684000
rect 4400 681000 526600 682600
rect 4400 679600 5400 681000
rect 7000 679600 9200 681000
rect 10800 679600 14000 681000
rect 15600 679600 526600 681000
rect 4400 678000 16600 679600
rect 4400 676600 5400 678000
rect 7000 676600 9200 678000
rect 10800 676600 14000 678000
rect 15600 676600 16600 678000
rect 4400 675000 16600 676600
rect 4400 673600 5400 675000
rect 7000 673600 9200 675000
rect 10800 673600 14000 675000
rect 15600 673600 16600 675000
rect 4400 672000 16600 673600
rect 4400 670600 5400 672000
rect 7000 670600 9200 672000
rect 10800 670600 14000 672000
rect 15600 670600 16600 672000
rect 4400 669000 16600 670600
rect 4400 667600 5400 669000
rect 7000 667600 9200 669000
rect 10800 667600 14000 669000
rect 15600 667600 16600 669000
rect 4400 666000 16600 667600
rect 4400 664600 5400 666000
rect 7000 664600 9200 666000
rect 10800 664600 14000 666000
rect 15600 664600 16600 666000
rect 4400 663000 16600 664600
rect 4400 661600 5400 663000
rect 7000 661600 9200 663000
rect 10800 661600 14000 663000
rect 15600 661600 16600 663000
rect 4400 660000 16600 661600
rect 4400 658600 5400 660000
rect 7000 658600 9200 660000
rect 10800 658600 14000 660000
rect 15600 658600 16600 660000
rect 4400 657000 16600 658600
rect 4400 655600 5400 657000
rect 7000 655600 9200 657000
rect 10800 655600 14000 657000
rect 15600 655600 16600 657000
rect 4400 654000 16600 655600
rect 4400 652600 5400 654000
rect 7000 652600 9200 654000
rect 10800 652600 14000 654000
rect 15600 652600 16600 654000
rect 4400 651000 16600 652600
rect 4400 649600 5400 651000
rect 7000 649600 9200 651000
rect 10800 649600 14000 651000
rect 15600 649600 16600 651000
rect -800 643842 1660 648642
rect 4400 648000 16600 649600
rect 4400 646600 5400 648000
rect 7000 646600 9200 648000
rect 10800 646600 14000 648000
rect 15600 646600 16600 648000
rect 4400 645000 16600 646600
rect 4400 643600 5400 645000
rect 7000 643600 9200 645000
rect 10800 643600 14000 645000
rect 15600 643600 16600 645000
rect 4400 642000 16600 643600
rect 4400 640600 5400 642000
rect 7000 640600 9200 642000
rect 10800 640600 14000 642000
rect 15600 640600 16600 642000
rect 4400 639000 16600 640600
rect -800 633842 1660 638642
rect 4400 637600 5400 639000
rect 7000 637600 9200 639000
rect 10800 637600 14000 639000
rect 15600 637600 16600 639000
rect 4400 636000 16600 637600
rect 4400 634600 5400 636000
rect 7000 634600 9200 636000
rect 10800 634600 14000 636000
rect 15600 634600 16600 636000
rect 4400 633000 16600 634600
rect 4400 631600 5400 633000
rect 7000 631600 9200 633000
rect 10800 631600 14000 633000
rect 15600 631600 16600 633000
rect 4400 630000 16600 631600
rect 4400 628600 5400 630000
rect 7000 628600 9200 630000
rect 10800 628600 14000 630000
rect 15600 628600 16600 630000
rect 4400 627000 16600 628600
rect 4400 625600 5400 627000
rect 7000 625600 9200 627000
rect 10800 625600 14000 627000
rect 15600 625600 16600 627000
rect 4400 624000 16600 625600
rect 4400 622600 5400 624000
rect 7000 622600 9200 624000
rect 10800 622600 14000 624000
rect 15600 622600 16600 624000
rect 4400 621000 16600 622600
rect 4400 619600 5400 621000
rect 7000 619600 9200 621000
rect 10800 619600 14000 621000
rect 15600 619600 16600 621000
rect 4400 618000 16600 619600
rect 4400 616600 5400 618000
rect 7000 616600 9200 618000
rect 10800 616600 14000 618000
rect 15600 616600 16600 618000
rect 4400 615000 16600 616600
rect 4400 613600 5400 615000
rect 7000 613600 9200 615000
rect 10800 613600 14000 615000
rect 15600 613600 16600 615000
rect 4400 612000 16600 613600
rect 4400 610600 5400 612000
rect 7000 610600 9200 612000
rect 10800 610600 14000 612000
rect 15600 610600 16600 612000
rect 4400 609000 16600 610600
rect 4400 607600 5400 609000
rect 7000 607600 9200 609000
rect 10800 607600 14000 609000
rect 15600 607600 16600 609000
rect 4400 606000 16600 607600
rect 4400 604600 5400 606000
rect 7000 604600 9200 606000
rect 10800 604600 14000 606000
rect 15600 604600 16600 606000
rect 4400 603000 16600 604600
rect 4400 601600 5400 603000
rect 7000 601600 9200 603000
rect 10800 601600 14000 603000
rect 15600 601600 16600 603000
rect 4400 600000 16600 601600
rect 4400 598600 5400 600000
rect 7000 598600 9200 600000
rect 10800 598600 14000 600000
rect 15600 598600 16600 600000
rect 4400 597000 16600 598600
rect 4400 595600 5400 597000
rect 7000 595600 9200 597000
rect 10800 595600 14000 597000
rect 15600 595600 16600 597000
rect 4400 594000 16600 595600
rect 4400 592600 5400 594000
rect 7000 592600 9200 594000
rect 10800 592600 14000 594000
rect 15600 592600 16600 594000
rect 4400 591000 16600 592600
rect 4400 589600 5400 591000
rect 7000 589600 9200 591000
rect 10800 589600 14000 591000
rect 15600 589600 16600 591000
rect 4400 588000 16600 589600
rect 4400 586600 5400 588000
rect 7000 586600 9200 588000
rect 10800 586600 14000 588000
rect 15600 586600 16600 588000
rect 4400 585000 16600 586600
rect 4400 583600 5400 585000
rect 7000 583600 9200 585000
rect 10800 583600 14000 585000
rect 15600 583600 16600 585000
rect 4400 582000 16600 583600
rect 4400 580600 5400 582000
rect 7000 580600 9200 582000
rect 10800 580600 14000 582000
rect 15600 580600 16600 582000
rect 4400 579000 16600 580600
rect 4400 577600 5400 579000
rect 7000 577600 9200 579000
rect 10800 577600 14000 579000
rect 15600 577600 16600 579000
rect 4400 576000 16600 577600
rect 4400 574600 5400 576000
rect 7000 574600 9200 576000
rect 10800 574600 14000 576000
rect 15600 574600 16600 576000
rect 4400 573000 16600 574600
rect 4400 571600 5400 573000
rect 7000 571600 9200 573000
rect 10800 571600 14000 573000
rect 15600 571600 16600 573000
rect 4400 570000 16600 571600
rect 4400 568600 5400 570000
rect 7000 568600 9200 570000
rect 10800 568600 14000 570000
rect 15600 568600 16600 570000
rect 4400 567000 16600 568600
rect 4400 565600 5400 567000
rect 7000 565600 9200 567000
rect 10800 565600 14000 567000
rect 15600 565600 16600 567000
rect 4400 564800 16600 565600
rect 475200 645200 477800 678200
rect 481200 677400 526600 679600
rect 580110 682990 583580 683510
rect 580110 678030 580470 682990
rect 581910 682984 583580 682990
rect 581910 678030 584800 682984
rect 580110 677984 584800 678030
rect 580110 677660 583580 677984
rect 481200 676200 494400 677400
rect 481200 674200 482800 676200
rect 493000 674200 494400 676200
rect 481200 673200 494400 674200
rect 481200 671200 482800 673200
rect 493000 671200 494400 673200
rect 481200 670200 494400 671200
rect 481200 668200 482800 670200
rect 493000 668200 494400 670200
rect 519680 669740 527080 670340
rect 481200 667200 494400 668200
rect 512600 668160 513720 668240
rect 512600 667690 512660 668160
rect 513650 667690 513720 668160
rect 512600 667610 513720 667690
rect 481200 665200 482800 667200
rect 493000 666000 494400 667200
rect 493000 665200 496400 666000
rect 481200 664200 496400 665200
rect 512350 665740 514050 667390
rect 512350 665220 514060 665740
rect 512350 664910 512420 665220
rect 514020 664910 514060 665220
rect 512350 664820 514060 664910
rect 519680 664340 520580 669740
rect 526480 664340 527080 669740
rect 481200 662200 482800 664200
rect 493000 662200 496400 664200
rect 481200 661200 496400 662200
rect 481200 659200 482800 661200
rect 493000 659200 496400 661200
rect 481200 658200 496400 659200
rect 481200 656200 482800 658200
rect 493000 656200 496400 658200
rect 481200 655200 496400 656200
rect 502600 664000 513200 664200
rect 502600 661000 505800 664000
rect 511400 661000 513200 664000
rect 519680 663640 527080 664340
rect 502600 660200 513200 661000
rect 502600 657200 505800 660200
rect 511400 659600 513200 660200
rect 511400 657200 516000 659600
rect 502600 656400 516000 657200
rect 502600 655600 509400 656400
rect 481200 653200 482800 655200
rect 493000 653800 496400 655200
rect 493000 653200 494400 653800
rect 508400 653600 509400 655600
rect 507200 653510 509400 653600
rect 481200 652200 494400 653200
rect 503450 653460 503690 653490
rect 503450 652270 503480 653460
rect 503670 652270 503690 653460
rect 503450 652240 503690 652270
rect 507070 653400 509400 653510
rect 515000 653400 516000 656400
rect 481200 650200 482800 652200
rect 493000 650200 494400 652200
rect 481200 649200 494400 650200
rect 481200 647200 482800 649200
rect 493000 647200 494400 649200
rect 481200 646200 494400 647200
rect 481200 645200 482800 646200
rect 475200 644200 482800 645200
rect 493000 644200 494400 646200
rect 475200 643200 494400 644200
rect 475200 641200 482800 643200
rect 493000 641200 494400 643200
rect 475200 640200 494400 641200
rect 475200 638200 482800 640200
rect 493000 638200 494400 640200
rect 475200 637200 494400 638200
rect 475200 635200 482800 637200
rect 493000 635200 494400 637200
rect 475200 634200 494400 635200
rect 475200 632200 482800 634200
rect 493000 632200 494400 634200
rect 475200 629800 494400 632200
rect 507070 650800 516000 653400
rect 507070 647800 509400 650800
rect 515000 647800 516000 650800
rect 507070 643400 516000 647800
rect 507070 640400 509400 643400
rect 515000 640400 516000 643400
rect 519780 646740 527180 647440
rect 519780 641340 520780 646740
rect 526680 641340 527180 646740
rect 519780 640740 527180 641340
rect 576350 644584 583900 644590
rect 576350 644270 584800 644584
rect 507070 637600 516000 640400
rect 507070 634600 509400 637600
rect 515000 634600 516000 637600
rect 507070 631810 516000 634600
rect 507200 631800 516000 631810
rect 507200 631200 509400 631800
rect 475200 570400 486400 629800
rect 508400 628800 509400 631200
rect 515000 628800 516000 631800
rect 576350 630020 576690 644270
rect 583530 639784 584800 644270
rect 583530 634584 583900 639784
rect 583530 630020 584800 634584
rect 576350 629784 584800 630020
rect 576350 629740 583900 629784
rect 508400 628200 516000 628800
rect 519880 623040 527180 623740
rect 519880 617740 520580 623040
rect 526580 617740 527180 623040
rect 519880 617040 527180 617740
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 497000 579200 503400 586200
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 577270 583674 583810 584240
rect 577270 583570 584800 583674
rect 577270 580390 577730 583570
rect 583180 583562 584800 583570
rect 583180 580390 583810 583562
rect 577270 579860 583810 580390
rect 1200 564730 17400 564800
rect 330 564400 17400 564730
rect 330 564320 4400 564400
rect 330 564242 870 564320
rect -800 559442 870 564242
rect 330 554242 870 559442
rect -800 549442 870 554242
rect 330 549250 870 549442
rect 2600 563000 4400 564320
rect 6000 563000 7200 564400
rect 8800 563000 9800 564400
rect 11400 563000 12800 564400
rect 14400 563000 15600 564400
rect 17200 563000 17400 564400
rect 2600 562200 15800 563000
rect 17000 562200 17400 563000
rect 2600 561600 17400 562200
rect 2600 561400 15800 561600
rect 17000 561400 17400 561600
rect 2600 560000 4400 561400
rect 6000 560000 7200 561400
rect 8800 560000 9800 561400
rect 11400 560000 12800 561400
rect 14400 560000 15600 561400
rect 17200 560000 17400 561400
rect 2600 559400 17400 560000
rect 2600 558200 15800 559400
rect 17000 558200 17400 559400
rect 2600 556800 4400 558200
rect 6000 556800 7200 558200
rect 8800 556800 9800 558200
rect 11400 556800 12800 558200
rect 14400 556800 15600 558200
rect 17200 556800 17400 558200
rect 2600 555800 15800 556800
rect 17000 555800 17400 556800
rect 2600 554400 4400 555800
rect 6000 554400 7200 555800
rect 8800 554400 9800 555800
rect 11400 554400 12800 555800
rect 14400 554400 15600 555800
rect 17200 554400 17400 555800
rect 2600 553400 15800 554400
rect 17000 553400 17400 554400
rect 2600 553200 17400 553400
rect 2600 551800 4400 553200
rect 6000 551800 7200 553200
rect 8800 551800 9800 553200
rect 11400 551800 12800 553200
rect 14400 551800 15600 553200
rect 17200 551800 17400 553200
rect 2600 551200 15800 551800
rect 17000 551200 17400 551800
rect 2600 550600 17400 551200
rect 2600 549250 4400 550600
rect 330 549200 4400 549250
rect 6000 549200 7200 550600
rect 8800 549200 9800 550600
rect 11400 549200 12800 550600
rect 14400 549200 15600 550600
rect 17200 549200 17400 550600
rect 330 548800 15800 549200
rect 17000 548800 17400 549200
rect 330 548720 16000 548800
rect 1200 548600 16000 548720
rect 16600 548600 17400 548800
rect 1200 548400 17400 548600
rect 475200 557400 488400 570400
rect 497000 568600 503200 579200
rect 511690 574080 519090 574680
rect 504810 572500 505930 572580
rect 504810 572030 504870 572500
rect 505860 572030 505930 572500
rect 504810 571950 505930 572030
rect 504560 570080 506260 571730
rect 504560 569560 506270 570080
rect 504560 569250 504630 569560
rect 506230 569250 506270 569560
rect 504560 569160 506270 569250
rect 494600 567600 503200 568600
rect 511690 568680 512590 574080
rect 518490 568680 519090 574080
rect 564280 574210 571680 574810
rect 557400 572630 558520 572710
rect 511690 567980 519090 568680
rect 529400 571400 539000 572400
rect 557400 572160 557460 572630
rect 558450 572160 558520 572630
rect 557400 572080 558520 572160
rect 494600 564600 497200 567600
rect 502800 566600 503200 567600
rect 502800 564600 508000 566600
rect 494600 563000 508000 564600
rect 494600 560000 501400 563000
rect 507000 560000 508000 563000
rect 494600 559800 508000 560000
rect 495460 557800 495700 557830
rect 6880 536700 7340 536740
rect 6880 534720 6920 536700
rect 7200 534720 7340 536700
rect 6880 534680 7340 534720
rect 8380 536700 8740 536740
rect 8380 534720 8420 536700
rect 8700 534720 8740 536700
rect 8380 534680 8740 534720
rect 475200 533800 486400 557400
rect 495460 556610 495490 557800
rect 495680 556610 495700 557800
rect 495460 556580 495700 556610
rect 499080 557800 499790 557850
rect 500400 557800 508000 559800
rect 499080 557400 508000 557800
rect 499080 554400 501400 557400
rect 507000 554400 508000 557400
rect 499080 550000 508000 554400
rect 529400 558400 541000 571400
rect 557150 569690 558860 571700
rect 557150 569380 557220 569690
rect 558820 569380 558860 569690
rect 557150 569290 558860 569380
rect 564280 568810 565180 574210
rect 571080 568810 571680 574210
rect 547200 567600 555800 568600
rect 564280 568110 571680 568810
rect 547200 564600 549800 567600
rect 555400 566800 555800 567600
rect 555400 564600 560400 566800
rect 547200 563600 560400 564600
rect 547200 560600 553800 563600
rect 559400 560600 560400 563600
rect 547200 560000 560400 560600
rect 552800 558400 560400 560000
rect 529400 554200 539000 558400
rect 551800 558000 560400 558400
rect 551800 557980 553800 558000
rect 548050 557930 548290 557960
rect 548050 556740 548080 557930
rect 548270 556740 548290 557930
rect 548050 556710 548290 556740
rect 499080 547000 501400 550000
rect 507000 547000 508000 550000
rect 499080 544200 508000 547000
rect 511790 551080 519190 551780
rect 511790 545680 512790 551080
rect 518690 545680 519190 551080
rect 511790 545080 519190 545680
rect 499080 541200 501400 544200
rect 507000 541200 508000 544200
rect 499080 538400 508000 541200
rect 499080 536150 501400 538400
rect 499400 535400 501400 536150
rect 507000 535400 508000 538400
rect 499400 535000 508000 535400
rect 500400 534800 508000 535000
rect 3230 532080 6770 532400
rect 3230 531700 3710 532080
rect 4140 531700 4930 532080
rect 5360 531700 6770 532080
rect 3230 531120 6770 531700
rect 3230 530740 3700 531120
rect 4130 530740 4920 531120
rect 5350 530740 6770 531120
rect 3230 530170 6770 530740
rect 3230 529790 3660 530170
rect 4090 529790 4880 530170
rect 5310 529790 6770 530170
rect 3230 529050 6770 529790
rect 3230 528670 3700 529050
rect 4130 528670 4920 529050
rect 5350 528670 6770 529050
rect 3230 528180 6770 528670
rect 3230 527800 3680 528180
rect 4110 527800 4900 528180
rect 5330 527800 6770 528180
rect 3230 527440 6770 527800
rect 475200 516200 485800 533800
rect 527800 533600 539000 554200
rect 551670 555000 553800 557980
rect 559400 555000 560400 558000
rect 551670 550600 560400 555000
rect 551670 547600 553800 550600
rect 559400 547600 560400 550600
rect 551670 544800 560400 547600
rect 564380 551210 571780 551910
rect 564380 545810 565380 551210
rect 571280 545810 571780 551210
rect 582340 550562 584800 555362
rect 564380 545210 571780 545810
rect 551670 541800 553800 544800
rect 559400 541800 560400 544800
rect 551670 540200 560400 541800
rect 582340 540562 584800 545362
rect 575600 540200 582600 540400
rect 551670 539000 582600 540200
rect 551670 536280 553800 539000
rect 551800 536000 553800 536280
rect 559400 536000 582600 539000
rect 551800 535200 582600 536000
rect 511890 527380 519190 528080
rect 511890 522080 512590 527380
rect 518590 522080 519190 527380
rect 511890 521380 519190 522080
rect 527800 516200 537400 533600
rect 557800 533200 582600 535200
rect 564480 527510 571780 528210
rect 564480 522210 565180 527510
rect 571180 522210 571780 527510
rect 564480 521510 571780 522210
rect 475200 515400 537400 516200
rect 160 512460 2530 512620
rect 160 511670 300 512460
rect 130 511642 300 511670
rect -800 511530 300 511642
rect 160 511100 300 511530
rect 2350 511100 2530 512460
rect 160 510950 2530 511100
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect 475200 506600 567600 515400
rect 575600 515200 582600 533200
rect -800 505620 480 505732
rect 190 469210 2560 469370
rect 190 468420 330 469210
rect -800 468308 330 468420
rect 190 467850 330 468308
rect 2380 467850 2560 469210
rect 190 467700 2560 467850
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect 1200 424800 10600 425100
rect 200 424600 10600 424800
rect 200 424016 400 424600
rect -800 423904 400 424016
rect 200 423400 400 423904
rect 1800 423400 10600 424600
rect 200 423200 10600 423400
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect 200 381300 2000 381500
rect 200 380794 400 381300
rect -800 380682 400 380794
rect 200 380100 400 380682
rect 1800 380100 2000 381300
rect 200 379900 2000 380100
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 600 375400 2400 375600
rect 600 375000 1000 375400
rect 2000 375000 2400 375400
rect 600 374800 2400 375000
rect 600 374400 1000 374800
rect 2000 374400 2400 374800
rect 600 374000 2400 374400
rect 600 373600 1000 374000
rect 2000 373600 2400 374000
rect 600 373200 2400 373600
rect 600 372800 1000 373200
rect 2000 372800 2400 373200
rect 600 372400 2400 372800
rect 600 372000 1000 372400
rect 2000 372000 2400 372400
rect 600 371600 2400 372000
rect 600 371200 1000 371600
rect 2000 371200 2400 371600
rect 600 370800 2400 371200
rect 600 370400 1000 370800
rect 2000 370400 2400 370800
rect 600 369400 2400 370400
rect 600 368800 800 369400
rect 1400 368800 2400 369400
rect 600 367400 2400 368800
rect 3200 368200 10600 423200
rect 600 366800 800 367400
rect 1400 366800 2400 367400
rect 2500 368000 10600 368200
rect 2500 367200 2700 368000
rect 10400 367200 10600 368000
rect 2500 367000 10600 367200
rect 15400 367100 17400 367300
rect 600 365400 2400 366800
rect 600 364800 800 365400
rect 1400 365140 2400 365400
rect 15400 366800 15800 367100
rect 17100 366800 17400 367100
rect 15400 366100 17400 366800
rect 15400 365800 15800 366100
rect 17100 365800 17400 366100
rect 1400 364800 2723 365140
rect 600 363400 2723 364800
rect 600 362800 800 363400
rect 1400 362800 2723 363400
rect 600 361400 2723 362800
rect 600 360800 800 361400
rect 1400 360800 2723 361400
rect 600 359400 2723 360800
rect 600 358800 800 359400
rect 1400 358800 2723 359400
rect 600 357400 2723 358800
rect 600 356800 800 357400
rect 1400 356800 2723 357400
rect 600 355400 2723 356800
rect 600 354800 800 355400
rect 1400 354800 2723 355400
rect 600 353400 2723 354800
rect 600 352800 800 353400
rect 1400 352800 2723 353400
rect 600 351400 2723 352800
rect 600 350800 800 351400
rect 1400 350800 2723 351400
rect 600 349400 2723 350800
rect 600 348800 800 349400
rect 1400 348800 2723 349400
rect 600 347400 2723 348800
rect 600 346800 800 347400
rect 1400 346800 2723 347400
rect 600 345400 2723 346800
rect 600 344800 800 345400
rect 1400 344800 2723 345400
rect 600 343440 2723 344800
rect 15400 365100 17400 365800
rect 15400 364800 15800 365100
rect 17100 364800 17400 365100
rect 15400 364100 17400 364800
rect 15400 363800 15800 364100
rect 17100 363800 17400 364100
rect 15400 363100 17400 363800
rect 15400 362800 15800 363100
rect 17100 362800 17400 363100
rect 15400 362100 17400 362800
rect 15400 361800 15800 362100
rect 17100 361800 17400 362100
rect 15400 361100 17400 361800
rect 15400 360800 15800 361100
rect 17100 360800 17400 361100
rect 15400 360100 17400 360800
rect 15400 359800 15800 360100
rect 17100 359800 17400 360100
rect 15400 359100 17400 359800
rect 15400 358800 15800 359100
rect 17100 358800 17400 359100
rect 15400 358100 17400 358800
rect 15400 357800 15800 358100
rect 17100 357800 17400 358100
rect 15400 357100 17400 357800
rect 15400 356800 15800 357100
rect 17100 356800 17400 357100
rect 15400 356100 17400 356800
rect 15400 355800 15800 356100
rect 17100 355800 17400 356100
rect 15400 355100 17400 355800
rect 15400 354800 15800 355100
rect 17100 354800 17400 355100
rect 15400 354100 17400 354800
rect 15400 353800 15800 354100
rect 17100 353800 17400 354100
rect 15400 353100 17400 353800
rect 15400 352800 15800 353100
rect 17100 352800 17400 353100
rect 15400 352100 17400 352800
rect 15400 351800 15800 352100
rect 17100 351800 17400 352100
rect 15400 351100 17400 351800
rect 15400 350800 15800 351100
rect 17100 350800 17400 351100
rect 15400 350100 17400 350800
rect 15400 349800 15800 350100
rect 17100 349800 17400 350100
rect 15400 349100 17400 349800
rect 15400 348800 15800 349100
rect 17100 348800 17400 349100
rect 15400 348100 17400 348800
rect 15400 347800 15800 348100
rect 17100 347800 17400 348100
rect 15400 347100 17400 347800
rect 15400 346800 15800 347100
rect 17100 346800 17400 347100
rect 15400 346100 17400 346800
rect 15400 345800 15800 346100
rect 17100 345800 17400 346100
rect 15400 345100 17400 345800
rect 15400 344800 15800 345100
rect 17100 344800 17400 345100
rect 6103 344680 6343 344710
rect 6103 343490 6123 344680
rect 6313 343490 6343 344680
rect 15400 344100 17400 344800
rect 15400 343800 15800 344100
rect 17100 343800 17400 344100
rect 15400 343700 17400 343800
rect 6103 343460 6343 343490
rect 600 341000 2400 343440
rect 600 339200 7200 341000
rect -800 338642 -187 338754
rect 200 338100 2000 338300
rect -800 337460 -187 337572
rect 200 336900 400 338100
rect 1800 336900 2000 338100
rect 200 336700 2000 336900
rect -800 336278 -187 336390
rect -800 335096 -187 335208
rect -800 333914 -187 334026
rect 2400 333200 7200 339200
rect 12700 340600 15400 341100
rect 12700 340300 13800 340600
rect 15000 340300 15400 340600
rect 12700 339600 15400 340300
rect 12700 339300 13800 339600
rect 15000 339300 15400 339600
rect 12700 338600 15400 339300
rect 12700 338300 13800 338600
rect 15000 338300 15400 338600
rect 12700 337600 15400 338300
rect 12700 337300 13800 337600
rect 15000 337300 15400 337600
rect 12700 336600 15400 337300
rect 12700 336300 13800 336600
rect 15000 336300 15400 336600
rect 12700 335600 15400 336300
rect 12700 335300 13800 335600
rect 15000 335300 15400 335600
rect 12700 334600 15400 335300
rect 12700 334300 13800 334600
rect 15000 334300 15400 334600
rect 12700 333600 15400 334300
rect 12700 333300 13800 333600
rect 15000 333300 15400 333600
rect 12700 333000 15400 333300
rect -800 332732 -187 332844
rect 2840 326413 5250 326483
rect 2840 324813 2930 326413
rect 3240 324813 5250 326413
rect 5630 326173 6260 326233
rect 5630 325183 5710 326173
rect 6180 325183 6260 326173
rect 5630 325113 6260 325183
rect 2840 324773 5250 324813
rect 200 296100 2000 296300
rect 200 295532 400 296100
rect -800 295420 400 295532
rect 200 294900 400 295420
rect 1800 294900 2000 296100
rect 200 294700 2000 294900
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 200 253000 2000 253200
rect 200 252510 400 253000
rect -800 252398 400 252510
rect 200 251800 400 252398
rect 1800 251800 2000 253000
rect 200 251600 2000 251800
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 400 177688 2740 177720
rect -800 177370 2740 177688
rect -800 172888 700 177370
rect 400 167688 700 172888
rect -800 163110 700 167688
rect 2330 163110 2740 177370
rect -800 162888 2740 163110
rect 400 162870 2740 162888
rect 200 125500 2000 125700
rect 200 124888 400 125500
rect -800 124776 400 124888
rect 200 124300 400 124776
rect 1800 124300 2000 125500
rect 200 124100 2000 124300
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect -800 16910 480 17022
rect -800 15728 480 15840
rect -800 14546 480 14658
rect -800 13364 480 13476
rect -800 12182 480 12294
rect -800 11000 480 11112
rect -800 9818 480 9930
rect -800 8636 480 8748
rect -800 7454 480 7566
rect -800 6272 480 6384
rect -800 5090 480 5202
rect -800 3908 480 4020
rect -800 2726 480 2838
rect 475200 2000 477800 506600
rect 530400 505800 567600 506600
rect 554600 503800 567600 505800
rect 571200 504800 582600 515200
rect 553290 496610 554540 496640
rect 553290 496420 553320 496610
rect 554510 496420 554540 496610
rect 553290 496400 554540 496420
rect 556800 494600 565200 497600
rect 571200 494600 578200 504800
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 556800 494400 578200 494600
rect 556800 494200 562000 494400
rect 532860 492800 554560 493020
rect 532400 491600 554600 492800
rect 556800 491600 557800 494200
rect 528400 490600 557800 491600
rect 528400 485000 529000 490600
rect 532000 485000 534800 490600
rect 537800 485000 540600 490600
rect 543600 485000 548000 490600
rect 551000 485000 553600 490600
rect 556600 488600 557800 490600
rect 560800 488800 562000 494200
rect 565000 492400 578200 494400
rect 580300 495690 582680 496130
rect 580300 493390 580590 495690
rect 582340 494930 582680 495690
rect 583520 495322 584800 495434
rect 582340 494252 583840 494930
rect 582340 494140 584800 494252
rect 582340 493400 583840 494140
rect 582340 493390 582680 493400
rect 580300 493190 582680 493390
rect 565000 488800 577000 492400
rect 560800 488600 577000 488800
rect 556600 488000 571000 488600
rect 556600 485000 559800 488000
rect 565870 487470 568440 487540
rect 565870 485870 565960 487470
rect 566270 485870 568440 487470
rect 568660 487230 569290 487290
rect 568660 486240 568740 487230
rect 569210 486240 569290 487230
rect 568660 486170 569290 486240
rect 565870 485840 568440 485870
rect 565870 485830 566790 485840
rect 528400 484000 559800 485000
rect 518090 479510 524790 480210
rect 518090 473510 518790 479510
rect 524090 473510 524790 479510
rect 518090 472910 524790 473510
rect 541790 479310 548490 480310
rect 541790 473410 542390 479310
rect 547790 473410 548490 479310
rect 541790 472910 548490 473410
rect 564690 479510 571390 480410
rect 564690 473610 565390 479510
rect 570790 473610 571390 479510
rect 564690 473010 571390 473610
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 576460 450970 578840 451410
rect 576460 448670 576750 450970
rect 578500 450600 578840 450970
rect 583520 450900 584800 451012
rect 578500 450540 583070 450600
rect 578500 449830 583860 450540
rect 578500 449718 584800 449830
rect 578500 448970 583860 449718
rect 578500 448880 583070 448970
rect 578500 448670 578840 448880
rect 576460 448470 578840 448670
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 571350 407140 583800 407350
rect 571350 405820 571720 407140
rect 577750 406590 583800 407140
rect 577750 406478 584800 406590
rect 577750 405820 583800 406478
rect 571350 405610 583800 405820
rect 583520 405296 584800 405408
rect 575600 365000 576200 365200
rect 578400 365000 579000 365200
rect 573800 364800 574800 365000
rect 573800 363400 574000 364800
rect 574600 363400 574800 364800
rect 573800 363200 574800 363400
rect 575600 363400 575800 365000
rect 576000 363400 576200 365000
rect 575600 363200 576200 363400
rect 576600 364800 577600 365000
rect 576600 363400 576800 364800
rect 577400 363400 577600 364800
rect 576600 363200 577600 363400
rect 578400 363400 578600 365000
rect 578800 363400 579000 365000
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 578400 363200 579000 363400
rect 583520 362420 584800 362532
rect 572400 361400 574800 361800
rect 572400 361200 572600 361400
rect 573400 361200 573800 361400
rect 574600 361200 574800 361400
rect 583520 361238 584800 361350
rect 572400 361000 574800 361200
rect 572400 360800 572600 361000
rect 573400 360800 573800 361000
rect 574600 360800 574800 361000
rect 572400 360600 574800 360800
rect 572400 360400 572600 360600
rect 573400 360400 573800 360600
rect 574600 360400 574800 360600
rect 572400 360200 574800 360400
rect 572400 360000 572600 360200
rect 573400 360000 573800 360200
rect 574600 360000 574800 360200
rect 572400 359800 574800 360000
rect 572400 359600 572600 359800
rect 573400 359600 573800 359800
rect 574600 359600 574800 359800
rect 572400 359400 574800 359600
rect 572400 359200 572600 359400
rect 573400 359200 573800 359400
rect 574600 359200 574800 359400
rect 579020 360800 583790 360900
rect 579020 359440 579150 360800
rect 582190 360168 583790 360800
rect 582190 360056 584800 360168
rect 582190 359440 583790 360056
rect 579020 359300 583790 359440
rect 572400 359000 574800 359200
rect 572400 358800 572600 359000
rect 573400 358800 573800 359000
rect 574600 358800 574800 359000
rect 583520 358874 584800 358986
rect 572400 358600 574800 358800
rect 572400 358400 572600 358600
rect 573400 358400 573800 358600
rect 574600 358400 574800 358600
rect 572400 358200 574800 358400
rect 572400 358000 572600 358200
rect 573400 358000 573800 358200
rect 574600 358000 574800 358200
rect 572400 357800 574800 358000
rect 572400 357600 572600 357800
rect 573400 357600 573800 357800
rect 574600 357600 574800 357800
rect 572400 357400 574800 357600
rect 572400 357200 572600 357400
rect 573400 357200 573800 357400
rect 574600 357200 574800 357400
rect 572400 357000 574800 357200
rect 572400 356800 572600 357000
rect 573400 356800 573800 357000
rect 574600 356800 574800 357000
rect 572400 356600 574800 356800
rect 572400 356400 572600 356600
rect 573400 356400 573800 356600
rect 574600 356400 574800 356600
rect 572400 356200 574800 356400
rect 572400 356000 572600 356200
rect 573400 356000 573800 356200
rect 574600 356000 574800 356200
rect 572400 355800 574800 356000
rect 572400 355600 572600 355800
rect 573400 355600 573800 355800
rect 574600 355600 574800 355800
rect 572400 355400 574800 355600
rect 572400 355200 572600 355400
rect 573400 355200 573800 355400
rect 574600 355200 574800 355400
rect 572400 355000 574800 355200
rect 572400 354800 572600 355000
rect 573400 354800 573800 355000
rect 574600 354800 574800 355000
rect 572400 354600 574800 354800
rect 572400 354400 572600 354600
rect 573400 354400 573800 354600
rect 574600 354400 574800 354600
rect 572400 354200 574800 354400
rect 572400 354000 572600 354200
rect 573400 354000 573800 354200
rect 574600 354000 574800 354200
rect 572400 353800 574800 354000
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 576850 315490 583800 315640
rect 576850 314100 576980 315490
rect 579620 314946 583800 315490
rect 579620 314834 584800 314946
rect 579620 314100 583800 314834
rect 576850 313990 583800 314100
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 566800 271600 572000 272000
rect 566800 270600 569200 271600
rect 571600 270600 572000 271600
rect 583520 271594 584800 271706
rect 566800 269600 572000 270600
rect 573510 270990 583830 271200
rect 573510 269790 573690 270990
rect 579290 270524 583830 270990
rect 579290 270412 584800 270524
rect 579290 269790 583830 270412
rect 573510 269620 583830 269790
rect 566800 268600 569200 269600
rect 571600 268600 572000 269600
rect 583520 269230 584800 269342
rect 566800 267600 572000 268600
rect 566800 266600 569200 267600
rect 571600 266600 572000 267600
rect 566800 265600 572000 266600
rect 566800 264600 569200 265600
rect 571600 264600 572000 265600
rect 566800 263600 572000 264600
rect 566800 262600 569200 263600
rect 571600 262600 572000 263600
rect 566800 261600 572000 262600
rect 566800 260600 569200 261600
rect 571600 260600 572000 261600
rect 566800 259600 572000 260600
rect 566800 258600 569200 259600
rect 571600 258600 572000 259600
rect 566800 258200 572000 258600
rect 580430 265330 583850 266510
rect 580430 264550 580810 265330
rect 583470 264550 583850 265330
rect 580430 263500 583850 264550
rect 580430 262720 580840 263500
rect 583500 262720 583850 263500
rect 580430 261910 583850 262720
rect 580430 261130 580810 261910
rect 583470 261130 583850 261910
rect 580430 260290 583850 261130
rect 580430 259510 580780 260290
rect 583440 259510 583850 260290
rect 580430 259100 583850 259510
rect 580430 258320 580810 259100
rect 583470 258320 583850 259100
rect 566800 241530 569360 258200
rect 580430 257890 583850 258320
rect 566800 241440 569770 241530
rect 566800 240400 569360 241440
rect 581280 241180 583800 257890
rect 581270 240910 583800 241180
rect 581270 240640 583750 240910
rect 581270 240400 581990 240640
rect 566800 238070 568630 240400
rect 566800 216370 568640 238070
rect 581250 224390 581990 240400
rect 572020 217610 572260 217640
rect 572020 216420 572040 217610
rect 572230 216420 572260 217610
rect 581250 217000 583800 224390
rect 572020 216390 572260 216420
rect 566800 216140 568310 216370
rect 566800 215720 568380 216140
rect 566850 213950 568380 215720
rect 566850 206040 574230 213950
rect 566850 205960 568380 206040
rect 580300 203600 583800 217000
rect 579200 201000 581200 201200
rect 579200 198160 579460 201000
rect 580960 198160 581200 201000
rect 579200 189900 579500 198160
rect 580900 189900 581200 198160
rect 579200 189500 581200 189900
rect 582300 196230 583800 203600
rect 582300 191430 584800 196230
rect 582300 186230 583800 191430
rect 582300 181430 584800 186230
rect 576200 175500 579600 175800
rect 576200 167200 576400 175500
rect 579400 167200 579600 175500
rect 576200 166600 579600 167200
rect 572900 152000 576700 152600
rect 572900 151830 573200 152000
rect 572900 148990 573150 151830
rect 572900 143700 573200 148990
rect 576200 143700 576700 152000
rect 572900 143300 576700 143700
rect 582300 151630 583800 181430
rect 582300 146830 584800 151630
rect 582300 141630 583800 146830
rect 582300 137300 584800 141630
rect 582340 136830 584800 137300
rect 570290 130870 578040 131480
rect 570290 130820 570900 130870
rect 570290 130770 570880 130820
rect 570290 123400 570850 130770
rect 577350 123400 578040 130870
rect 570290 123020 578040 123400
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 583520 13364 584800 13476
rect 583520 12182 584800 12294
rect 583520 11000 584800 11112
rect 583520 9818 584800 9930
rect 583520 8636 584800 8748
rect 583520 7454 584800 7566
rect 583520 6272 584800 6384
rect 583520 5090 584800 5202
rect 583520 3908 584800 4020
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 228670 701850 232530 702520
rect 222600 698000 226600 698800
rect 222600 696800 226600 697600
rect 222600 695600 226600 696400
rect 330480 701740 334340 702410
rect 324200 698000 328200 698800
rect 324200 696800 328200 697600
rect 324200 695600 328200 696400
rect 510880 696600 525130 703440
rect 482800 674200 493000 676200
rect 482800 671200 493000 673200
rect 482800 668200 493000 670200
rect 512660 667690 513650 668160
rect 482800 665200 493000 667200
rect 520580 664340 526480 669740
rect 482800 662200 493000 664200
rect 482800 659200 493000 661200
rect 482800 656200 493000 658200
rect 505800 661000 511400 664000
rect 505800 657200 511400 660200
rect 482800 653200 493000 655200
rect 503480 652270 503670 653460
rect 509400 653400 515000 656400
rect 482800 650200 493000 652200
rect 482800 647200 493000 649200
rect 482800 644200 493000 646200
rect 482800 641200 493000 643200
rect 482800 638200 493000 640200
rect 482800 635200 493000 637200
rect 482800 632200 493000 634200
rect 509400 647800 515000 650800
rect 509400 640400 515000 643400
rect 520780 641340 526680 646740
rect 509400 634600 515000 637600
rect 509400 628800 515000 631800
rect 576690 630020 583530 644270
rect 520580 617740 526580 623040
rect 870 549250 2600 564320
rect 15800 563000 17000 563600
rect 15800 562200 17000 563000
rect 15800 561400 17000 561600
rect 15800 560200 17000 561400
rect 15800 558200 17000 559400
rect 15800 558000 17000 558200
rect 15800 556800 17000 557200
rect 15800 555800 17000 556800
rect 15800 554400 17000 554800
rect 15800 553400 17000 554400
rect 15800 551800 17000 552600
rect 15800 551600 16000 551800
rect 16000 551600 16600 551800
rect 16600 551600 17000 551800
rect 15800 551200 17000 551600
rect 15800 549200 17000 550200
rect 15800 548800 16000 549200
rect 16000 548800 16600 549200
rect 16600 548800 17000 549200
rect 504870 572030 505860 572500
rect 512590 568680 518490 574080
rect 557460 572160 558450 572630
rect 497200 564600 502800 567600
rect 501400 560000 507000 563000
rect 6920 534720 7200 536700
rect 8420 534720 8700 536700
rect 495490 556610 495680 557800
rect 501400 554400 507000 557400
rect 565180 568810 571080 574210
rect 549800 564600 555400 567600
rect 553800 560600 559400 563600
rect 548080 556740 548270 557930
rect 501400 547000 507000 550000
rect 512790 545680 518690 551080
rect 501400 541200 507000 544200
rect 501400 535400 507000 538400
rect 3710 531700 4140 532080
rect 4930 531700 5360 532080
rect 3700 530740 4130 531120
rect 4920 530740 5350 531120
rect 3660 529790 4090 530170
rect 4880 529790 5310 530170
rect 3700 528670 4130 529050
rect 4920 528670 5350 529050
rect 3680 527800 4110 528180
rect 4900 527800 5330 528180
rect 553800 555000 559400 558000
rect 553800 547600 559400 550600
rect 565380 545810 571280 551210
rect 553800 541800 559400 544800
rect 553800 536000 559400 539000
rect 512590 522080 518590 527380
rect 565180 522210 571180 527510
rect 1000 375000 2000 375400
rect 1000 374400 2000 374800
rect 1000 373600 2000 374000
rect 1000 372800 2000 373200
rect 1000 372000 2000 372400
rect 1000 371200 2000 371600
rect 1000 370400 2000 370800
rect 800 368800 1400 369400
rect 800 366800 1400 367400
rect 2700 367200 10400 368000
rect 800 364800 1400 365400
rect 15800 366800 17100 367100
rect 15800 365800 17100 366100
rect 800 362800 1400 363400
rect 800 360800 1400 361400
rect 800 358800 1400 359400
rect 800 356800 1400 357400
rect 800 354800 1400 355400
rect 800 352800 1400 353400
rect 800 350800 1400 351400
rect 800 348800 1400 349400
rect 800 346800 1400 347400
rect 800 344800 1400 345400
rect 15800 364800 17100 365100
rect 15800 363800 17100 364100
rect 15800 362800 17100 363100
rect 15800 361800 17100 362100
rect 15800 360800 17100 361100
rect 15800 359800 17100 360100
rect 15800 358800 17100 359100
rect 15800 357800 17100 358100
rect 15800 356800 17100 357100
rect 15800 355800 17100 356100
rect 15800 354800 17100 355100
rect 15800 353800 17100 354100
rect 15800 352800 17100 353100
rect 15800 351800 17100 352100
rect 15800 350800 17100 351100
rect 15800 349800 17100 350100
rect 15800 348800 17100 349100
rect 15800 347800 17100 348100
rect 15800 346800 17100 347100
rect 15800 345800 17100 346100
rect 15800 344800 17100 345100
rect 6123 343490 6313 344680
rect 15800 343800 17100 344100
rect 13800 340300 15000 340600
rect 13800 339300 15000 339600
rect 13800 338300 15000 338600
rect 13800 337300 15000 337600
rect 13800 336300 15000 336600
rect 13800 335300 15000 335600
rect 13800 334300 15000 334600
rect 13800 333300 15000 333600
rect 5710 325183 6180 326173
rect 700 163110 2330 177370
rect 553320 496420 554510 496610
rect 529000 485000 532000 490600
rect 534800 485000 537800 490600
rect 540600 485000 543600 490600
rect 548000 485000 551000 490600
rect 553600 485000 556600 490600
rect 557800 488600 560800 494200
rect 562000 488800 565000 494400
rect 568740 486240 569210 487230
rect 518790 473510 524090 479510
rect 542390 473410 547790 479310
rect 565390 473610 570790 479510
rect 574000 363400 574600 364800
rect 575800 363400 576000 365000
rect 576800 363400 577400 364800
rect 578600 363400 578800 365000
rect 572600 361200 573400 361400
rect 573800 361200 574600 361400
rect 572600 360800 573400 361000
rect 573800 360800 574600 361000
rect 572600 360400 573400 360600
rect 573800 360400 574600 360600
rect 572600 360000 573400 360200
rect 573800 360000 574600 360200
rect 572600 359600 573400 359800
rect 573800 359600 574600 359800
rect 572600 359200 573400 359400
rect 573800 359200 574600 359400
rect 572600 358800 573400 359000
rect 573800 358800 574600 359000
rect 572600 358400 573400 358600
rect 573800 358400 574600 358600
rect 572600 358000 573400 358200
rect 573800 358000 574600 358200
rect 572600 357600 573400 357800
rect 573800 357600 574600 357800
rect 572600 357200 573400 357400
rect 573800 357200 574600 357400
rect 572600 356800 573400 357000
rect 573800 356800 574600 357000
rect 572600 356400 573400 356600
rect 573800 356400 574600 356600
rect 572600 356000 573400 356200
rect 573800 356000 574600 356200
rect 572600 355600 573400 355800
rect 573800 355600 574600 355800
rect 572600 355200 573400 355400
rect 573800 355200 574600 355400
rect 572600 354800 573400 355000
rect 573800 354800 574600 355000
rect 572600 354400 573400 354600
rect 573800 354400 574600 354600
rect 572600 354000 573400 354200
rect 573800 354000 574600 354200
rect 569200 270600 571600 271600
rect 569200 268600 571600 269600
rect 569200 266600 571600 267600
rect 569200 264600 571600 265600
rect 569200 262600 571600 263600
rect 569200 260600 571600 261600
rect 569200 258600 571600 259600
rect 580810 264550 583470 265330
rect 580840 262720 583500 263500
rect 580810 261130 583470 261910
rect 580780 259510 583440 260290
rect 580810 258320 583470 259100
rect 572040 216420 572230 217610
rect 579460 198160 580960 201000
rect 579500 189900 580900 198160
rect 576400 167200 579400 175500
rect 573200 151830 576200 152000
rect 573150 148990 576200 151830
rect 573200 143700 576200 148990
rect 570900 130820 577350 130870
rect 570900 123430 577350 130820
<< mimcap >>
rect 512450 667010 513950 667290
rect 512450 666100 512730 667010
rect 513640 666100 513950 667010
rect 512450 665790 513950 666100
rect 504660 571350 506160 571630
rect 504660 570440 504940 571350
rect 505850 570440 506160 571350
rect 557590 571230 558220 571290
rect 557590 570740 557670 571230
rect 558130 570740 558220 571230
rect 557590 570660 558220 570740
rect 504660 570130 506160 570440
rect 566840 487160 568340 487440
rect 566840 486250 567150 487160
rect 568060 486250 568340 487160
rect 566840 485940 568340 486250
rect 4210 325963 4840 326043
rect 4210 325503 4290 325963
rect 4780 325503 4840 325963
rect 4210 325413 4840 325503
<< mimcapcontact >>
rect 512730 666100 513640 667010
rect 504940 570440 505850 571350
rect 557670 570740 558130 571230
rect 567150 486250 568060 487160
rect 4290 325503 4780 325963
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702990 232594 704800
rect 227594 702520 233090 702990
rect 227594 702300 228670 702520
rect 228240 701850 228670 702300
rect 232530 701850 233090 702520
rect 318994 702300 323994 704800
rect 329294 702880 334294 704800
rect 510600 703440 525450 703780
rect 329294 702410 334900 702880
rect 329294 702300 330480 702410
rect 228240 701380 233090 701850
rect 330050 701740 330480 702300
rect 334340 701740 334900 702410
rect 330050 701270 334900 701740
rect 222200 698800 227200 699600
rect 222200 698000 222600 698800
rect 226600 698000 227200 698800
rect 222200 697600 227200 698000
rect 222200 696800 222600 697600
rect 226600 696800 227200 697600
rect 222200 696400 227200 696800
rect 222200 695600 222600 696400
rect 226600 695600 227200 696400
rect 222200 695400 227200 695600
rect 323800 698800 328800 699600
rect 323800 698000 324200 698800
rect 328200 698000 328800 698800
rect 323800 697600 328800 698000
rect 323800 696800 324200 697600
rect 328200 696800 328800 697600
rect 323800 696400 328800 696800
rect 323800 695600 324200 696400
rect 328200 695600 328800 696400
rect 510600 696600 510880 703440
rect 525130 696600 525450 703440
rect 510600 696230 525450 696600
rect 510600 696200 525400 696230
rect 323800 695400 328800 695600
rect 222200 694400 227200 695000
rect 535200 694600 555000 695200
rect 524200 694400 566600 694600
rect 3800 691800 566600 694400
rect 3800 691600 535600 691800
rect 3800 690200 7200 691600
rect 9000 690200 11000 691600
rect 12800 691400 535600 691600
rect 12800 690200 15800 691400
rect 16800 690200 18800 691400
rect 19800 690200 21800 691400
rect 22800 690200 24800 691400
rect 25800 690200 27800 691400
rect 28800 690200 30800 691400
rect 31800 690200 33800 691400
rect 34800 690200 36800 691400
rect 37800 690200 39800 691400
rect 40800 690200 42800 691400
rect 43800 690200 45800 691400
rect 46800 690200 48800 691400
rect 49800 690200 51800 691400
rect 52800 690200 54800 691400
rect 55800 690200 57800 691400
rect 58800 690200 60800 691400
rect 61800 690200 63800 691400
rect 64800 690200 66800 691400
rect 67800 690200 69800 691400
rect 70800 690200 72800 691400
rect 73800 690200 75800 691400
rect 76800 690200 78800 691400
rect 79800 690200 81800 691400
rect 82800 690200 84800 691400
rect 85800 690200 87800 691400
rect 88800 690200 90800 691400
rect 91800 690200 93800 691400
rect 94800 690200 96800 691400
rect 97800 690200 99800 691400
rect 100800 690200 102800 691400
rect 103800 690200 105800 691400
rect 106800 690200 108800 691400
rect 109800 690200 111800 691400
rect 112800 690200 114800 691400
rect 115800 690200 117800 691400
rect 118800 690200 120800 691400
rect 121800 690200 123800 691400
rect 124800 690200 126800 691400
rect 127800 690200 129800 691400
rect 130800 690200 132800 691400
rect 133800 690200 135800 691400
rect 136800 690200 138800 691400
rect 139800 690200 141800 691400
rect 142800 690200 144800 691400
rect 145800 690200 147800 691400
rect 148800 690200 150800 691400
rect 151800 690200 153800 691400
rect 154800 690200 156800 691400
rect 157800 690200 159800 691400
rect 160800 690200 162800 691400
rect 163800 690200 165800 691400
rect 166800 690200 168800 691400
rect 169800 690200 171800 691400
rect 172800 690200 174800 691400
rect 175800 690200 177800 691400
rect 178800 690200 180800 691400
rect 181800 690200 183800 691400
rect 184800 690200 186800 691400
rect 187800 690200 189800 691400
rect 190800 690200 192800 691400
rect 193800 690200 195800 691400
rect 196800 690200 198800 691400
rect 199800 690200 201800 691400
rect 202800 690200 204800 691400
rect 205800 690200 207800 691400
rect 208800 690200 210800 691400
rect 211800 690200 213800 691400
rect 214800 690200 216800 691400
rect 217800 690200 219800 691400
rect 220800 690200 222800 691400
rect 223800 690200 225800 691400
rect 226800 690200 228800 691400
rect 229800 690200 231800 691400
rect 232800 690200 234800 691400
rect 235800 690200 237800 691400
rect 238800 690200 240800 691400
rect 241800 690200 243800 691400
rect 244800 690200 246800 691400
rect 247800 690200 249800 691400
rect 250800 690200 252800 691400
rect 253800 690200 255800 691400
rect 256800 690200 258800 691400
rect 259800 690200 261800 691400
rect 262800 690200 264800 691400
rect 265800 690200 267800 691400
rect 268800 690200 270800 691400
rect 271800 690200 273800 691400
rect 274800 690200 276800 691400
rect 277800 690200 279800 691400
rect 280800 690200 282800 691400
rect 283800 690200 285800 691400
rect 286800 690200 288800 691400
rect 289800 690200 291800 691400
rect 292800 690200 294800 691400
rect 295800 690200 297800 691400
rect 298800 690200 300800 691400
rect 301800 690200 303800 691400
rect 304800 690200 306800 691400
rect 307800 690200 309800 691400
rect 310800 690200 312800 691400
rect 313800 690200 315800 691400
rect 316800 690200 318800 691400
rect 319800 690200 321800 691400
rect 322800 690200 324800 691400
rect 325800 690200 327800 691400
rect 328800 690200 330800 691400
rect 331800 690200 333800 691400
rect 334800 690200 336800 691400
rect 337800 690200 339800 691400
rect 340800 690200 342800 691400
rect 343800 690200 345800 691400
rect 346800 690200 348800 691400
rect 349800 690200 351800 691400
rect 352800 690200 354800 691400
rect 355800 690200 357800 691400
rect 358800 690200 360800 691400
rect 361800 690200 363800 691400
rect 364800 690200 366800 691400
rect 367800 690200 369800 691400
rect 370800 690200 372800 691400
rect 373800 690200 375800 691400
rect 376800 690200 378800 691400
rect 379800 690200 381800 691400
rect 382800 690200 384800 691400
rect 385800 690200 387800 691400
rect 388800 690200 390800 691400
rect 391800 690200 393800 691400
rect 394800 690200 396800 691400
rect 397800 690200 399800 691400
rect 400800 690200 402800 691400
rect 403800 690200 405800 691400
rect 406800 690200 408800 691400
rect 409800 690200 411800 691400
rect 412800 690200 414800 691400
rect 415800 690200 417800 691400
rect 418800 690200 420800 691400
rect 421800 690200 423800 691400
rect 424800 690200 426800 691400
rect 427800 690200 429800 691400
rect 430800 690200 432800 691400
rect 433800 690200 435800 691400
rect 436800 690200 438800 691400
rect 439800 690200 441800 691400
rect 442800 690200 444800 691400
rect 445800 690200 447800 691400
rect 448800 690200 450800 691400
rect 451800 690200 453800 691400
rect 454800 690200 456800 691400
rect 457800 690200 459800 691400
rect 460800 690200 462800 691400
rect 463800 690200 465800 691400
rect 466800 690200 468800 691400
rect 469800 690200 471800 691400
rect 472800 690200 474800 691400
rect 475800 690200 477800 691400
rect 478800 690200 480800 691400
rect 481800 690200 483800 691400
rect 484800 690200 486800 691400
rect 487800 690200 489800 691400
rect 490800 690200 492800 691400
rect 493800 690200 495800 691400
rect 496800 690200 498800 691400
rect 499800 690200 501800 691400
rect 502800 690200 504800 691400
rect 505800 690200 507800 691400
rect 508800 690200 510800 691400
rect 511800 690200 513800 691400
rect 514800 690200 516800 691400
rect 517800 690200 519800 691400
rect 520800 690200 522800 691400
rect 523800 690200 525800 691400
rect 526800 690200 528800 691400
rect 529800 690200 531800 691400
rect 532800 690200 535600 691400
rect 3800 689800 535600 690200
rect 544200 689800 545600 691800
rect 554200 689800 566600 691800
rect 3800 688600 566600 689800
rect 3800 687200 7200 688600
rect 9000 687200 11000 688600
rect 12800 688400 566600 688600
rect 12800 687200 15800 688400
rect 16800 687200 18800 688400
rect 19800 687200 21800 688400
rect 22800 687200 24800 688400
rect 25800 687200 27800 688400
rect 28800 687200 30800 688400
rect 31800 687200 33800 688400
rect 34800 687200 36800 688400
rect 37800 687200 39800 688400
rect 40800 687200 42800 688400
rect 43800 687200 45800 688400
rect 46800 687200 48800 688400
rect 49800 687200 51800 688400
rect 52800 687200 54800 688400
rect 55800 687200 57800 688400
rect 58800 687200 60800 688400
rect 61800 687200 63800 688400
rect 64800 687200 66800 688400
rect 67800 687200 69800 688400
rect 70800 687200 72800 688400
rect 73800 687200 75800 688400
rect 76800 687200 78800 688400
rect 79800 687200 81800 688400
rect 82800 687200 84800 688400
rect 85800 687200 87800 688400
rect 88800 687200 90800 688400
rect 91800 687200 93800 688400
rect 94800 687200 96800 688400
rect 97800 687200 99800 688400
rect 100800 687200 102800 688400
rect 103800 687200 105800 688400
rect 106800 687200 108800 688400
rect 109800 687200 111800 688400
rect 112800 687200 114800 688400
rect 115800 687200 117800 688400
rect 118800 687200 120800 688400
rect 121800 687200 123800 688400
rect 124800 687200 126800 688400
rect 127800 687200 129800 688400
rect 130800 687200 132800 688400
rect 133800 687200 135800 688400
rect 136800 687200 138800 688400
rect 139800 687200 141800 688400
rect 142800 687200 144800 688400
rect 145800 687200 147800 688400
rect 148800 687200 150800 688400
rect 151800 687200 153800 688400
rect 154800 687200 156800 688400
rect 157800 687200 159800 688400
rect 160800 687200 162800 688400
rect 163800 687200 165800 688400
rect 166800 687200 168800 688400
rect 169800 687200 171800 688400
rect 172800 687200 174800 688400
rect 175800 687200 177800 688400
rect 178800 687200 180800 688400
rect 181800 687200 183800 688400
rect 184800 687200 186800 688400
rect 187800 687200 189800 688400
rect 190800 687200 192800 688400
rect 193800 687200 195800 688400
rect 196800 687200 198800 688400
rect 199800 687200 201800 688400
rect 202800 687200 204800 688400
rect 205800 687200 207800 688400
rect 208800 687200 210800 688400
rect 211800 687200 213800 688400
rect 214800 687200 216800 688400
rect 217800 687200 219800 688400
rect 220800 687200 222800 688400
rect 223800 687200 225800 688400
rect 226800 687200 228800 688400
rect 229800 687200 231800 688400
rect 232800 687200 234800 688400
rect 235800 687200 237800 688400
rect 238800 687200 240800 688400
rect 241800 687200 243800 688400
rect 244800 687200 246800 688400
rect 247800 687200 249800 688400
rect 250800 687200 252800 688400
rect 253800 687200 255800 688400
rect 256800 687200 258800 688400
rect 259800 687200 261800 688400
rect 262800 687200 264800 688400
rect 265800 687200 267800 688400
rect 268800 687200 270800 688400
rect 271800 687200 273800 688400
rect 274800 687200 276800 688400
rect 277800 687200 279800 688400
rect 280800 687200 282800 688400
rect 283800 687200 285800 688400
rect 286800 687200 288800 688400
rect 289800 687200 291800 688400
rect 292800 687200 294800 688400
rect 295800 687200 297800 688400
rect 298800 687200 300800 688400
rect 301800 687200 303800 688400
rect 304800 687200 306800 688400
rect 307800 687200 309800 688400
rect 310800 687200 312800 688400
rect 313800 687200 315800 688400
rect 316800 687200 318800 688400
rect 319800 687200 321800 688400
rect 322800 687200 324800 688400
rect 325800 687200 327800 688400
rect 328800 687200 330800 688400
rect 331800 687200 333800 688400
rect 334800 687200 336800 688400
rect 337800 687200 339800 688400
rect 340800 687200 342800 688400
rect 343800 687200 345800 688400
rect 346800 687200 348800 688400
rect 349800 687200 351800 688400
rect 352800 687200 354800 688400
rect 355800 687200 357800 688400
rect 358800 687200 360800 688400
rect 361800 687200 363800 688400
rect 364800 687200 366800 688400
rect 367800 687200 369800 688400
rect 370800 687200 372800 688400
rect 373800 687200 375800 688400
rect 376800 687200 378800 688400
rect 379800 687200 381800 688400
rect 382800 687200 384800 688400
rect 385800 687200 387800 688400
rect 388800 687200 390800 688400
rect 391800 687200 393800 688400
rect 394800 687200 396800 688400
rect 397800 687200 399800 688400
rect 400800 687200 402800 688400
rect 403800 687200 405800 688400
rect 406800 687200 408800 688400
rect 409800 687200 411800 688400
rect 412800 687200 414800 688400
rect 415800 687200 417800 688400
rect 418800 687200 420800 688400
rect 421800 687200 423800 688400
rect 424800 687200 426800 688400
rect 427800 687200 429800 688400
rect 430800 687200 432800 688400
rect 433800 687200 435800 688400
rect 436800 687200 438800 688400
rect 439800 687200 441800 688400
rect 442800 687200 444800 688400
rect 445800 687200 447800 688400
rect 448800 687200 450800 688400
rect 451800 687200 453800 688400
rect 454800 687200 456800 688400
rect 457800 687200 459800 688400
rect 460800 687200 462800 688400
rect 463800 687200 465800 688400
rect 466800 687200 468800 688400
rect 469800 687200 471800 688400
rect 472800 687200 474800 688400
rect 475800 687200 477800 688400
rect 478800 687200 480800 688400
rect 481800 687200 483800 688400
rect 484800 687200 486800 688400
rect 487800 687200 489800 688400
rect 490800 687200 492800 688400
rect 493800 687200 495800 688400
rect 496800 687200 498800 688400
rect 499800 687200 501800 688400
rect 502800 687200 504800 688400
rect 505800 687200 507800 688400
rect 508800 687200 510800 688400
rect 511800 687200 513800 688400
rect 514800 687200 516800 688400
rect 517800 687200 519800 688400
rect 520800 687200 522800 688400
rect 523800 687200 525800 688400
rect 526800 687200 528800 688400
rect 529800 687200 531800 688400
rect 532800 687800 566600 688400
rect 532800 687200 535600 687800
rect 3800 685800 535600 687200
rect 544200 685800 545600 687800
rect 554200 685800 566600 687800
rect 3800 685600 566600 685800
rect 3800 684200 7200 685600
rect 9000 684200 11000 685600
rect 12800 685400 566600 685600
rect 12800 684200 15800 685400
rect 16800 684200 18800 685400
rect 19800 684200 21800 685400
rect 22800 684200 24800 685400
rect 25800 684200 27800 685400
rect 28800 684200 30800 685400
rect 31800 684200 33800 685400
rect 34800 684200 36800 685400
rect 37800 684200 39800 685400
rect 40800 684200 42800 685400
rect 43800 684200 45800 685400
rect 46800 684200 48800 685400
rect 49800 684200 51800 685400
rect 52800 684200 54800 685400
rect 55800 684200 57800 685400
rect 58800 684200 60800 685400
rect 61800 684200 63800 685400
rect 64800 684200 66800 685400
rect 67800 684200 69800 685400
rect 70800 684200 72800 685400
rect 73800 684200 75800 685400
rect 76800 684200 78800 685400
rect 79800 684200 81800 685400
rect 82800 684200 84800 685400
rect 85800 684200 87800 685400
rect 88800 684200 90800 685400
rect 91800 684200 93800 685400
rect 94800 684200 96800 685400
rect 97800 684200 99800 685400
rect 100800 684200 102800 685400
rect 103800 684200 105800 685400
rect 106800 684200 108800 685400
rect 109800 684200 111800 685400
rect 112800 684200 114800 685400
rect 115800 684200 117800 685400
rect 118800 684200 120800 685400
rect 121800 684200 123800 685400
rect 124800 684200 126800 685400
rect 127800 684200 129800 685400
rect 130800 684200 132800 685400
rect 133800 684200 135800 685400
rect 136800 684200 138800 685400
rect 139800 684200 141800 685400
rect 142800 684200 144800 685400
rect 145800 684200 147800 685400
rect 148800 684200 150800 685400
rect 151800 684200 153800 685400
rect 154800 684200 156800 685400
rect 157800 684200 159800 685400
rect 160800 684200 162800 685400
rect 163800 684200 165800 685400
rect 166800 684200 168800 685400
rect 169800 684200 171800 685400
rect 172800 684200 174800 685400
rect 175800 684200 177800 685400
rect 178800 684200 180800 685400
rect 181800 684200 183800 685400
rect 184800 684200 186800 685400
rect 187800 684200 189800 685400
rect 190800 684200 192800 685400
rect 193800 684200 195800 685400
rect 196800 684200 198800 685400
rect 199800 684200 201800 685400
rect 202800 684200 204800 685400
rect 205800 684200 207800 685400
rect 208800 684200 210800 685400
rect 211800 684200 213800 685400
rect 214800 684200 216800 685400
rect 217800 684200 219800 685400
rect 220800 684200 222800 685400
rect 223800 684200 225800 685400
rect 226800 684200 228800 685400
rect 229800 684200 231800 685400
rect 232800 684200 234800 685400
rect 235800 684200 237800 685400
rect 238800 684200 240800 685400
rect 241800 684200 243800 685400
rect 244800 684200 246800 685400
rect 247800 684200 249800 685400
rect 250800 684200 252800 685400
rect 253800 684200 255800 685400
rect 256800 684200 258800 685400
rect 259800 684200 261800 685400
rect 262800 684200 264800 685400
rect 265800 684200 267800 685400
rect 268800 684200 270800 685400
rect 271800 684200 273800 685400
rect 274800 684200 276800 685400
rect 277800 684200 279800 685400
rect 280800 684200 282800 685400
rect 283800 684200 285800 685400
rect 286800 684200 288800 685400
rect 289800 684200 291800 685400
rect 292800 684200 294800 685400
rect 295800 684200 297800 685400
rect 298800 684200 300800 685400
rect 301800 684200 303800 685400
rect 304800 684200 306800 685400
rect 307800 684200 309800 685400
rect 310800 684200 312800 685400
rect 313800 684200 315800 685400
rect 316800 684200 318800 685400
rect 319800 684200 321800 685400
rect 322800 684200 324800 685400
rect 325800 684200 327800 685400
rect 328800 684200 330800 685400
rect 331800 684200 333800 685400
rect 334800 684200 336800 685400
rect 337800 684200 339800 685400
rect 340800 684200 342800 685400
rect 343800 684200 345800 685400
rect 346800 684200 348800 685400
rect 349800 684200 351800 685400
rect 352800 684200 354800 685400
rect 355800 684200 357800 685400
rect 358800 684200 360800 685400
rect 361800 684200 363800 685400
rect 364800 684200 366800 685400
rect 367800 684200 369800 685400
rect 370800 684200 372800 685400
rect 373800 684200 375800 685400
rect 376800 684200 378800 685400
rect 379800 684200 381800 685400
rect 382800 684200 384800 685400
rect 385800 684200 387800 685400
rect 388800 684200 390800 685400
rect 391800 684200 393800 685400
rect 394800 684200 396800 685400
rect 397800 684200 399800 685400
rect 400800 684200 402800 685400
rect 403800 684200 405800 685400
rect 406800 684200 408800 685400
rect 409800 684200 411800 685400
rect 412800 684200 414800 685400
rect 415800 684200 417800 685400
rect 418800 684200 420800 685400
rect 421800 684200 423800 685400
rect 424800 684200 426800 685400
rect 427800 684200 429800 685400
rect 430800 684200 432800 685400
rect 433800 684200 435800 685400
rect 436800 684200 438800 685400
rect 439800 684200 441800 685400
rect 442800 684200 444800 685400
rect 445800 684200 447800 685400
rect 448800 684200 450800 685400
rect 451800 684200 453800 685400
rect 454800 684200 456800 685400
rect 457800 684200 459800 685400
rect 460800 684200 462800 685400
rect 463800 684200 465800 685400
rect 466800 684200 468800 685400
rect 469800 684200 471800 685400
rect 472800 684200 474800 685400
rect 475800 684200 477800 685400
rect 478800 684200 480800 685400
rect 481800 684200 483800 685400
rect 484800 684200 486800 685400
rect 487800 684200 489800 685400
rect 490800 684200 492800 685400
rect 493800 684200 495800 685400
rect 496800 684200 498800 685400
rect 499800 684200 501800 685400
rect 502800 684200 504800 685400
rect 505800 684200 507800 685400
rect 508800 684200 510800 685400
rect 511800 684200 513800 685400
rect 514800 684200 516800 685400
rect 517800 684200 519800 685400
rect 520800 684200 522800 685400
rect 523800 684200 525800 685400
rect 526800 684200 528800 685400
rect 529800 684200 531800 685400
rect 532800 684200 566600 685400
rect 3800 683800 566600 684200
rect 3800 682600 535600 683800
rect 3800 681200 7200 682600
rect 9000 681200 11000 682600
rect 12800 682400 535600 682600
rect 12800 681200 15800 682400
rect 16800 681200 18800 682400
rect 19800 681200 21800 682400
rect 22800 681200 24800 682400
rect 25800 681200 27800 682400
rect 28800 681200 30800 682400
rect 31800 681200 33800 682400
rect 34800 681200 36800 682400
rect 37800 681200 39800 682400
rect 40800 681200 42800 682400
rect 43800 681200 45800 682400
rect 46800 681200 48800 682400
rect 49800 681200 51800 682400
rect 52800 681200 54800 682400
rect 55800 681200 57800 682400
rect 58800 681200 60800 682400
rect 61800 681200 63800 682400
rect 64800 681200 66800 682400
rect 67800 681200 69800 682400
rect 70800 681200 72800 682400
rect 73800 681200 75800 682400
rect 76800 681200 78800 682400
rect 79800 681200 81800 682400
rect 82800 681200 84800 682400
rect 85800 681200 87800 682400
rect 88800 681200 90800 682400
rect 91800 681200 93800 682400
rect 94800 681200 96800 682400
rect 97800 681200 99800 682400
rect 100800 681200 102800 682400
rect 103800 681200 105800 682400
rect 106800 681200 108800 682400
rect 109800 681200 111800 682400
rect 112800 681200 114800 682400
rect 115800 681200 117800 682400
rect 118800 681200 120800 682400
rect 121800 681200 123800 682400
rect 124800 681200 126800 682400
rect 127800 681200 129800 682400
rect 130800 681200 132800 682400
rect 133800 681200 135800 682400
rect 136800 681200 138800 682400
rect 139800 681200 141800 682400
rect 142800 681200 144800 682400
rect 145800 681200 147800 682400
rect 148800 681200 150800 682400
rect 151800 681200 153800 682400
rect 154800 681200 156800 682400
rect 157800 681200 159800 682400
rect 160800 681200 162800 682400
rect 163800 681200 165800 682400
rect 166800 681200 168800 682400
rect 169800 681200 171800 682400
rect 172800 681200 174800 682400
rect 175800 681200 177800 682400
rect 178800 681200 180800 682400
rect 181800 681200 183800 682400
rect 184800 681200 186800 682400
rect 187800 681200 189800 682400
rect 190800 681200 192800 682400
rect 193800 681200 195800 682400
rect 196800 681200 198800 682400
rect 199800 681200 201800 682400
rect 202800 681200 204800 682400
rect 205800 681200 207800 682400
rect 208800 681200 210800 682400
rect 211800 681200 213800 682400
rect 214800 681200 216800 682400
rect 217800 681200 219800 682400
rect 220800 681200 222800 682400
rect 223800 681200 225800 682400
rect 226800 681200 228800 682400
rect 229800 681200 231800 682400
rect 232800 681200 234800 682400
rect 235800 681200 237800 682400
rect 238800 681200 240800 682400
rect 241800 681200 243800 682400
rect 244800 681200 246800 682400
rect 247800 681200 249800 682400
rect 250800 681200 252800 682400
rect 253800 681200 255800 682400
rect 256800 681200 258800 682400
rect 259800 681200 261800 682400
rect 262800 681200 264800 682400
rect 265800 681200 267800 682400
rect 268800 681200 270800 682400
rect 271800 681200 273800 682400
rect 274800 681200 276800 682400
rect 277800 681200 279800 682400
rect 280800 681200 282800 682400
rect 283800 681200 285800 682400
rect 286800 681200 288800 682400
rect 289800 681200 291800 682400
rect 292800 681200 294800 682400
rect 295800 681200 297800 682400
rect 298800 681200 300800 682400
rect 301800 681200 303800 682400
rect 304800 681200 306800 682400
rect 307800 681200 309800 682400
rect 310800 681200 312800 682400
rect 313800 681200 315800 682400
rect 316800 681200 318800 682400
rect 319800 681200 321800 682400
rect 322800 681200 324800 682400
rect 325800 681200 327800 682400
rect 328800 681200 330800 682400
rect 331800 681200 333800 682400
rect 334800 681200 336800 682400
rect 337800 681200 339800 682400
rect 340800 681200 342800 682400
rect 343800 681200 345800 682400
rect 346800 681200 348800 682400
rect 349800 681200 351800 682400
rect 352800 681200 354800 682400
rect 355800 681200 357800 682400
rect 358800 681200 360800 682400
rect 361800 681200 363800 682400
rect 364800 681200 366800 682400
rect 367800 681200 369800 682400
rect 370800 681200 372800 682400
rect 373800 681200 375800 682400
rect 376800 681200 378800 682400
rect 379800 681200 381800 682400
rect 382800 681200 384800 682400
rect 385800 681200 387800 682400
rect 388800 681200 390800 682400
rect 391800 681200 393800 682400
rect 394800 681200 396800 682400
rect 397800 681200 399800 682400
rect 400800 681200 402800 682400
rect 403800 681200 405800 682400
rect 406800 681200 408800 682400
rect 409800 681200 411800 682400
rect 412800 681200 414800 682400
rect 415800 681200 417800 682400
rect 418800 681200 420800 682400
rect 421800 681200 423800 682400
rect 424800 681200 426800 682400
rect 427800 681200 429800 682400
rect 430800 681200 432800 682400
rect 433800 681200 435800 682400
rect 436800 681200 438800 682400
rect 439800 681200 441800 682400
rect 442800 681200 444800 682400
rect 445800 681200 447800 682400
rect 448800 681200 450800 682400
rect 451800 681200 453800 682400
rect 454800 681200 456800 682400
rect 457800 681200 459800 682400
rect 460800 681200 462800 682400
rect 463800 681200 465800 682400
rect 466800 681200 468800 682400
rect 469800 681200 471800 682400
rect 472800 681200 474800 682400
rect 475800 681200 477800 682400
rect 478800 681200 480800 682400
rect 481800 681200 483800 682400
rect 484800 681200 486800 682400
rect 487800 681200 489800 682400
rect 490800 681200 492800 682400
rect 493800 681200 495800 682400
rect 496800 681200 498800 682400
rect 499800 681200 501800 682400
rect 502800 681200 504800 682400
rect 505800 681200 507800 682400
rect 508800 681200 510800 682400
rect 511800 681200 513800 682400
rect 514800 681200 516800 682400
rect 517800 681200 519800 682400
rect 520800 681200 522800 682400
rect 523800 681200 525800 682400
rect 526800 681200 528800 682400
rect 529800 681200 531800 682400
rect 532800 681800 535600 682400
rect 544200 681800 545600 683800
rect 554200 681800 566600 683800
rect 532800 681200 566600 681800
rect 3800 679800 566600 681200
rect 3800 679600 535600 679800
rect 3800 678200 7200 679600
rect 9000 678200 11000 679600
rect 12800 678200 15000 679600
rect 3800 676600 15000 678200
rect 3800 675200 7200 676600
rect 9000 675200 11000 676600
rect 12800 675200 15000 676600
rect 3800 673600 15000 675200
rect 3800 672200 7200 673600
rect 9000 672200 11000 673600
rect 12800 672200 15000 673600
rect 3800 670600 15000 672200
rect 3800 669200 7200 670600
rect 9000 669200 11000 670600
rect 12800 669200 15000 670600
rect 3800 667600 15000 669200
rect 3800 666200 7200 667600
rect 9000 666200 11000 667600
rect 12800 666200 15000 667600
rect 3800 664600 15000 666200
rect 3800 663200 7200 664600
rect 9000 663200 11000 664600
rect 12800 663200 15000 664600
rect 3800 661600 15000 663200
rect 3800 660200 7200 661600
rect 9000 660200 11000 661600
rect 12800 660200 15000 661600
rect 3800 658600 15000 660200
rect 3800 657200 7200 658600
rect 9000 657200 11000 658600
rect 12800 657200 15000 658600
rect 3800 656000 15000 657200
rect 3800 654800 4800 656000
rect 6200 655600 15000 656000
rect 6200 654800 7200 655600
rect 3800 654200 7200 654800
rect 9000 654200 11000 655600
rect 12800 654200 15000 655600
rect 3800 654000 15000 654200
rect 3800 653800 4800 654000
rect 600 652800 4800 653800
rect 6200 652800 15000 654000
rect 600 652600 15000 652800
rect 600 652000 7200 652600
rect 600 650800 4800 652000
rect 6200 651200 7200 652000
rect 9000 651200 11000 652600
rect 12800 651200 15000 652600
rect 6200 650800 15000 651200
rect 600 650000 15000 650800
rect 600 648800 4800 650000
rect 6200 649600 15000 650000
rect 6200 648800 7200 649600
rect 600 648200 7200 648800
rect 9000 648200 11000 649600
rect 12800 648200 15000 649600
rect 600 648000 15000 648200
rect 600 646800 4800 648000
rect 6200 646800 15000 648000
rect 600 646600 15000 646800
rect 600 646000 7200 646600
rect 600 644800 4800 646000
rect 6200 645200 7200 646000
rect 9000 645200 11000 646600
rect 12800 645200 15000 646600
rect 6200 644800 15000 645200
rect 600 644000 15000 644800
rect 600 642800 4800 644000
rect 6200 643600 15000 644000
rect 6200 642800 7200 643600
rect 600 642200 7200 642800
rect 9000 642200 11000 643600
rect 12800 642200 15000 643600
rect 600 642000 15000 642200
rect 600 640800 4800 642000
rect 6200 640800 15000 642000
rect 600 640600 15000 640800
rect 600 640000 7200 640600
rect 600 638800 4800 640000
rect 6200 639200 7200 640000
rect 9000 639200 11000 640600
rect 12800 639200 15000 640600
rect 6200 638800 15000 639200
rect 600 638000 15000 638800
rect 600 636800 4800 638000
rect 6200 637600 15000 638000
rect 6200 636800 7200 637600
rect 600 636200 7200 636800
rect 9000 636200 11000 637600
rect 12800 636200 15000 637600
rect 600 636000 15000 636200
rect 600 634800 4800 636000
rect 6200 634800 15000 636000
rect 600 634600 15000 634800
rect 600 634000 7200 634600
rect 600 632800 4800 634000
rect 6200 633200 7200 634000
rect 9000 633200 11000 634600
rect 12800 633200 15000 634600
rect 6200 632800 15000 633200
rect 600 632000 15000 632800
rect 600 631800 4800 632000
rect 4400 630800 4800 631800
rect 6200 630800 7400 632000
rect 8800 631800 15000 632000
rect 475200 677400 477800 678200
rect 475200 676000 475800 677400
rect 477200 676000 477800 677400
rect 534800 677800 535600 679600
rect 544200 677800 545600 679800
rect 554200 679600 566600 679800
rect 554200 677800 555400 679600
rect 475200 675400 477800 676000
rect 475200 674000 475800 675400
rect 477200 674000 477800 675400
rect 475200 673400 477800 674000
rect 475200 672000 475800 673400
rect 477200 672000 477800 673400
rect 475200 671400 477800 672000
rect 475200 670000 475800 671400
rect 477200 670000 477800 671400
rect 475200 669400 477800 670000
rect 475200 668000 475800 669400
rect 477200 668000 477800 669400
rect 475200 667400 477800 668000
rect 475200 666000 475800 667400
rect 477200 666000 477800 667400
rect 475200 665400 477800 666000
rect 475200 664000 475800 665400
rect 477200 664000 477800 665400
rect 475200 663400 477800 664000
rect 475200 662000 475800 663400
rect 477200 662000 477800 663400
rect 475200 661400 477800 662000
rect 475200 660000 475800 661400
rect 477200 660000 477800 661400
rect 475200 659400 477800 660000
rect 475200 658000 475800 659400
rect 477200 658000 477800 659400
rect 475200 657400 477800 658000
rect 475200 656000 475800 657400
rect 477200 656000 477800 657400
rect 475200 655400 477800 656000
rect 475200 654000 475800 655400
rect 477200 654000 477800 655400
rect 475200 653400 477800 654000
rect 475200 652000 475800 653400
rect 477200 652000 477800 653400
rect 475200 651400 477800 652000
rect 475200 650000 475800 651400
rect 477200 650000 477800 651400
rect 475200 649400 477800 650000
rect 475200 648000 475800 649400
rect 477200 648000 477800 649400
rect 475200 647400 477800 648000
rect 475200 646000 475800 647400
rect 477200 646000 477800 647400
rect 475200 645400 477800 646000
rect 475200 644000 475800 645400
rect 477200 645200 477800 645400
rect 481200 676200 494400 677000
rect 481200 674200 482800 676200
rect 493000 674200 494400 676200
rect 481200 673200 494400 674200
rect 481200 671200 482800 673200
rect 493000 671200 494400 673200
rect 481200 670200 494400 671200
rect 534800 675800 555400 677800
rect 534800 673800 535600 675800
rect 544200 673800 545600 675800
rect 554200 673800 555400 675800
rect 534800 671800 555400 673800
rect 481200 668200 482800 670200
rect 493000 668200 494400 670200
rect 519680 669740 527080 670340
rect 481200 667200 494400 668200
rect 481200 665200 482800 667200
rect 493000 666000 494400 667200
rect 512600 668160 513720 668240
rect 512600 667690 512660 668160
rect 513650 667690 513720 668160
rect 512600 667010 513720 667690
rect 512600 666100 512730 667010
rect 513640 666100 513720 667010
rect 512600 666020 513720 666100
rect 493000 665200 496400 666000
rect 481200 664200 496400 665200
rect 519680 664340 520580 669740
rect 526480 664340 527080 669740
rect 481200 662200 482800 664200
rect 493000 662200 496400 664200
rect 481200 661200 496400 662200
rect 481200 659200 482800 661200
rect 493000 659200 496400 661200
rect 481200 658200 496400 659200
rect 481200 656200 482800 658200
rect 493000 656200 496400 658200
rect 481200 655200 496400 656200
rect 504600 664000 513200 664200
rect 504600 661000 505800 664000
rect 511400 661000 513200 664000
rect 519680 663640 527080 664340
rect 534800 669800 535600 671800
rect 544200 669800 545600 671800
rect 554200 669800 555400 671800
rect 534800 667800 555400 669800
rect 534800 665800 535600 667800
rect 544200 665800 545600 667800
rect 554200 665800 555400 667800
rect 534800 663800 555400 665800
rect 504600 660200 513200 661000
rect 504600 657200 505800 660200
rect 511400 659600 513200 660200
rect 534800 661800 535600 663800
rect 544200 661800 545600 663800
rect 554200 661800 555400 663800
rect 534800 659800 555400 661800
rect 511400 657200 516000 659600
rect 504600 656400 516000 657200
rect 504600 655600 509400 656400
rect 481200 653200 482800 655200
rect 493000 653800 496400 655200
rect 493000 653200 494400 653800
rect 481200 652200 494400 653200
rect 503450 653460 503690 653490
rect 503450 652270 503480 653460
rect 503670 653060 503690 653460
rect 508400 653400 509400 655600
rect 515000 653400 516000 656400
rect 503670 652660 507780 653060
rect 503670 652270 503690 652660
rect 503450 652240 503690 652270
rect 481200 650200 482800 652200
rect 493000 650200 494400 652200
rect 481200 649200 494400 650200
rect 481200 647200 482800 649200
rect 493000 647200 494400 649200
rect 481200 646200 494400 647200
rect 481200 645200 482800 646200
rect 477200 644200 482800 645200
rect 493000 644200 494400 646200
rect 477200 644000 494400 644200
rect 475200 643400 494400 644000
rect 475200 642000 475800 643400
rect 477200 643200 494400 643400
rect 477200 642000 482800 643200
rect 475200 641400 482800 642000
rect 475200 640000 475800 641400
rect 477200 641200 482800 641400
rect 493000 641200 494400 643200
rect 477200 640200 494400 641200
rect 477200 640000 482800 640200
rect 475200 639400 482800 640000
rect 475200 638000 475800 639400
rect 477200 638200 482800 639400
rect 493000 638200 494400 640200
rect 477200 638000 494400 638200
rect 475200 637400 494400 638000
rect 475200 636000 475800 637400
rect 477200 637200 494400 637400
rect 477200 636000 482800 637200
rect 475200 635400 482800 636000
rect 475200 634000 475800 635400
rect 477200 635200 482800 635400
rect 493000 635200 494400 637200
rect 477200 634200 494400 635200
rect 477200 634000 482800 634200
rect 475200 633400 482800 634000
rect 475200 632000 475800 633400
rect 477200 632200 482800 633400
rect 493000 632200 494400 634200
rect 477200 632000 494400 632200
rect 8800 630800 9200 631800
rect 4400 630000 9200 630800
rect 475200 631400 494400 632000
rect 4400 628800 4800 630000
rect 6200 628800 7400 630000
rect 8800 628800 9200 630000
rect 4400 628000 9200 628800
rect 4400 626800 4800 628000
rect 6200 626800 7400 628000
rect 8800 626800 9200 628000
rect 4400 626000 9200 626800
rect 4400 624800 4800 626000
rect 6200 624800 7400 626000
rect 8800 624800 9200 626000
rect 4400 624000 9200 624800
rect 4400 622800 4800 624000
rect 6200 622800 7400 624000
rect 8800 622800 9200 624000
rect 4400 622000 9200 622800
rect 4400 620800 4800 622000
rect 6200 620800 7400 622000
rect 8800 620800 9200 622000
rect 4400 620000 9200 620800
rect 4400 618800 4800 620000
rect 6200 618800 7400 620000
rect 8800 618800 9200 620000
rect 4400 618000 9200 618800
rect 4400 616800 4800 618000
rect 6200 616800 7400 618000
rect 8800 616800 9200 618000
rect 4400 616000 9200 616800
rect 4400 614800 4800 616000
rect 6200 614800 7400 616000
rect 8800 614800 9200 616000
rect 4400 614000 9200 614800
rect 4400 612800 4800 614000
rect 6200 612800 7400 614000
rect 8800 612800 9200 614000
rect 4400 612000 9200 612800
rect 4400 610800 4800 612000
rect 6200 610800 7400 612000
rect 8800 610800 9200 612000
rect 4400 610000 9200 610800
rect 4400 608800 4800 610000
rect 6200 608800 7400 610000
rect 8800 608800 9200 610000
rect 4400 608000 9200 608800
rect 4400 606800 4800 608000
rect 6200 606800 7400 608000
rect 8800 606800 9200 608000
rect 4400 606000 9200 606800
rect 4400 604800 4800 606000
rect 6200 604800 7400 606000
rect 8800 604800 9200 606000
rect 4400 604000 9200 604800
rect 4400 602800 4800 604000
rect 6200 602800 7400 604000
rect 8800 602800 9200 604000
rect 4400 602000 9200 602800
rect 4400 600800 4800 602000
rect 6200 600800 7400 602000
rect 8800 600800 9200 602000
rect 4400 600000 9200 600800
rect 4400 598800 4800 600000
rect 6200 598800 7400 600000
rect 8800 598800 9200 600000
rect 4400 598000 9200 598800
rect 4400 596800 4800 598000
rect 6200 596800 7400 598000
rect 8800 596800 9200 598000
rect 4400 596000 9200 596800
rect 4400 594800 4800 596000
rect 6200 594800 7400 596000
rect 8800 594800 9200 596000
rect 4400 594000 9200 594800
rect 4400 592800 4800 594000
rect 6200 592800 7400 594000
rect 8800 592800 9200 594000
rect 4400 592000 9200 592800
rect 4400 590800 4800 592000
rect 6200 590800 7400 592000
rect 8800 590800 9200 592000
rect 4400 590000 9200 590800
rect 4400 588800 4800 590000
rect 6200 588800 7400 590000
rect 8800 588800 9200 590000
rect 4400 588000 9200 588800
rect 4400 586800 4800 588000
rect 6200 586800 7400 588000
rect 8800 586800 9200 588000
rect 4400 586000 9200 586800
rect 4400 584800 4800 586000
rect 6200 584800 7400 586000
rect 8800 584800 9200 586000
rect 4400 584000 9200 584800
rect 4400 582800 4800 584000
rect 6200 582800 7400 584000
rect 8800 582800 9200 584000
rect 4400 582000 9200 582800
rect 4400 580800 4800 582000
rect 6200 580800 7400 582000
rect 8800 580800 9200 582000
rect 4400 580000 9200 580800
rect 4400 578800 4800 580000
rect 6200 578800 7400 580000
rect 8800 578800 9200 580000
rect 4400 578000 9200 578800
rect 4400 576800 4800 578000
rect 6200 576800 7400 578000
rect 8800 576800 9200 578000
rect 4400 576000 9200 576800
rect 4400 574800 4800 576000
rect 6200 574800 7400 576000
rect 8800 574800 9200 576000
rect 4400 574000 9200 574800
rect 4400 572800 4800 574000
rect 6200 572800 7400 574000
rect 8800 572800 9200 574000
rect 4400 572000 9200 572800
rect 4400 570800 4800 572000
rect 6200 570800 7400 572000
rect 8800 570800 9200 572000
rect 4400 570000 9200 570800
rect 4400 568800 4800 570000
rect 6200 568800 7400 570000
rect 8800 568800 9200 570000
rect 4400 568000 9200 568800
rect 4400 566800 4800 568000
rect 6200 566800 7400 568000
rect 8800 566800 9200 568000
rect 4400 566000 9200 566800
rect 4400 564800 4800 566000
rect 6200 564800 7400 566000
rect 8800 564800 9200 566000
rect 330 564320 2800 564730
rect 330 549250 870 564320
rect 2600 549250 2800 564320
rect 330 548720 2800 549250
rect 2700 548600 2800 548720
rect 4400 564000 9200 564800
rect 15800 630200 17000 630400
rect 15800 629600 16000 630200
rect 16800 629600 17000 630200
rect 15800 627200 17000 629600
rect 15800 626600 16000 627200
rect 16800 626600 17000 627200
rect 15800 624200 17000 626600
rect 15800 623600 16000 624200
rect 16800 623600 17000 624200
rect 15800 621200 17000 623600
rect 15800 620600 16000 621200
rect 16800 620600 17000 621200
rect 15800 618200 17000 620600
rect 15800 617600 16000 618200
rect 16800 617600 17000 618200
rect 15800 615200 17000 617600
rect 15800 614600 16000 615200
rect 16800 614600 17000 615200
rect 15800 612200 17000 614600
rect 15800 611600 16000 612200
rect 16800 611600 17000 612200
rect 15800 609200 17000 611600
rect 15800 608600 16000 609200
rect 16800 608600 17000 609200
rect 15800 606200 17000 608600
rect 15800 605600 16000 606200
rect 16800 605600 17000 606200
rect 15800 603200 17000 605600
rect 15800 602600 16000 603200
rect 16800 602600 17000 603200
rect 15800 600200 17000 602600
rect 15800 599600 16000 600200
rect 16800 599600 17000 600200
rect 15800 597200 17000 599600
rect 15800 596600 16000 597200
rect 16800 596600 17000 597200
rect 15800 594200 17000 596600
rect 15800 593600 16000 594200
rect 16800 593600 17000 594200
rect 15800 591200 17000 593600
rect 15800 590600 16000 591200
rect 16800 590600 17000 591200
rect 15800 588200 17000 590600
rect 15800 587600 16000 588200
rect 16800 587600 17000 588200
rect 15800 585200 17000 587600
rect 15800 584600 16000 585200
rect 16800 584600 17000 585200
rect 15800 582200 17000 584600
rect 15800 581600 16000 582200
rect 16800 581600 17000 582200
rect 15800 579200 17000 581600
rect 15800 578600 16000 579200
rect 16800 578600 17000 579200
rect 15800 576200 17000 578600
rect 15800 575600 16000 576200
rect 16800 575600 17000 576200
rect 15800 573200 17000 575600
rect 15800 572600 16000 573200
rect 16800 572600 17000 573200
rect 15800 570200 17000 572600
rect 15800 569600 16000 570200
rect 16800 569600 17000 570200
rect 15800 567200 17000 569600
rect 15800 566600 16000 567200
rect 16800 566600 17000 567200
rect 15800 564700 17000 566600
rect 475200 630000 475800 631400
rect 477200 630000 494400 631400
rect 475200 629800 494400 630000
rect 507660 629960 507780 652660
rect 503210 629880 507780 629960
rect 475200 629400 486400 629800
rect 475200 628000 475800 629400
rect 477200 628000 486400 629400
rect 475200 627400 486400 628000
rect 475200 626000 475800 627400
rect 477200 626000 486400 627400
rect 499220 629570 507780 629880
rect 508400 650800 516000 653400
rect 508400 647800 509400 650800
rect 515000 647800 516000 650800
rect 508400 643400 516000 647800
rect 534800 657800 535600 659800
rect 544200 657800 545600 659800
rect 554200 657800 555400 659800
rect 534800 655800 555400 657800
rect 534800 653800 535600 655800
rect 544200 653800 545600 655800
rect 554200 653800 555400 655800
rect 534800 651800 555400 653800
rect 534800 649800 535600 651800
rect 544200 649800 545600 651800
rect 554200 649800 555400 651800
rect 534800 647800 555400 649800
rect 508400 640400 509400 643400
rect 515000 640400 516000 643400
rect 519780 646740 527180 647440
rect 519780 641340 520780 646740
rect 526680 641340 527180 646740
rect 519780 640740 527180 641340
rect 534800 645800 535600 647800
rect 544200 645800 545600 647800
rect 554200 645800 555400 647800
rect 534800 643800 555400 645800
rect 534800 641800 535600 643800
rect 544200 641800 545600 643800
rect 554200 641800 555400 643800
rect 534800 641600 555400 641800
rect 556200 641600 566600 679600
rect 576350 644270 583900 644590
rect 576350 641600 576690 644270
rect 508400 637600 516000 640400
rect 508400 634600 509400 637600
rect 515000 635600 516000 637600
rect 534800 639800 576690 641600
rect 534800 637800 535600 639800
rect 544200 637800 545600 639800
rect 554200 637800 576690 639800
rect 534800 635800 576690 637800
rect 534800 635600 535600 635800
rect 515000 634600 535600 635600
rect 508400 633800 535600 634600
rect 544200 633800 545600 635800
rect 554200 633800 576690 635800
rect 508400 632000 576690 633800
rect 508400 631800 566600 632000
rect 499220 629510 507100 629570
rect 499220 628360 499340 629510
rect 507010 628360 507100 629510
rect 499220 627120 507100 628360
rect 508400 628800 509400 631800
rect 515000 629800 535600 631800
rect 544200 629800 545600 631800
rect 554200 629800 566600 631800
rect 515000 629000 566600 629800
rect 576350 630020 576690 632000
rect 583530 630020 583900 644270
rect 576350 629740 583900 630020
rect 515000 628800 561400 629000
rect 508400 628600 561400 628800
rect 508400 628200 516000 628600
rect 475200 625400 486400 626000
rect 475200 624000 475800 625400
rect 477200 624000 486400 625400
rect 475200 623400 486400 624000
rect 475200 622000 475800 623400
rect 477200 622000 486400 623400
rect 475200 621400 486400 622000
rect 475200 620000 475800 621400
rect 477200 620000 486400 621400
rect 475200 619400 486400 620000
rect 475200 618000 475800 619400
rect 477200 618000 486400 619400
rect 475200 617400 486400 618000
rect 475200 616000 475800 617400
rect 477200 616000 486400 617400
rect 519880 623040 527180 623740
rect 519880 617740 520580 623040
rect 526580 617740 527180 623040
rect 519880 617040 527180 617740
rect 475200 615400 486400 616000
rect 475200 614000 475800 615400
rect 477200 614000 486400 615400
rect 475200 613400 486400 614000
rect 475200 612000 475800 613400
rect 477200 612000 486400 613400
rect 475200 611400 486400 612000
rect 475200 610000 475800 611400
rect 477200 610000 486400 611400
rect 475200 609400 486400 610000
rect 475200 608000 475800 609400
rect 477200 608000 486400 609400
rect 475200 607400 486400 608000
rect 475200 606000 475800 607400
rect 477200 606000 486400 607400
rect 475200 605400 486400 606000
rect 475200 604000 475800 605400
rect 477200 604000 486400 605400
rect 475200 603400 486400 604000
rect 475200 602000 475800 603400
rect 477200 602000 486400 603400
rect 475200 601400 486400 602000
rect 475200 600000 475800 601400
rect 477200 600000 486400 601400
rect 551800 601200 561400 628600
rect 475200 599400 486400 600000
rect 475200 598000 475800 599400
rect 477200 598000 486400 599400
rect 475200 597400 486400 598000
rect 475200 596000 475800 597400
rect 477200 596000 486400 597400
rect 475200 595400 486400 596000
rect 475200 594000 475800 595400
rect 477200 594000 486400 595400
rect 549600 594400 561400 601200
rect 475200 593400 486400 594000
rect 475200 592000 475800 593400
rect 477200 592000 486400 593400
rect 475200 591400 486400 592000
rect 475200 590000 475800 591400
rect 477200 590000 486400 591400
rect 475200 589400 486400 590000
rect 475200 588000 475800 589400
rect 477200 588000 486400 589400
rect 475200 587400 486400 588000
rect 475200 586000 475800 587400
rect 477200 586000 486400 587400
rect 475200 585400 486400 586000
rect 475200 584000 475800 585400
rect 477200 584000 486400 585400
rect 475200 583400 486400 584000
rect 475200 582000 475800 583400
rect 477200 582000 486400 583400
rect 475200 581400 486400 582000
rect 475200 580000 475800 581400
rect 477200 580000 486400 581400
rect 475200 579400 486400 580000
rect 475200 578000 475800 579400
rect 477200 578000 486400 579400
rect 475200 577400 486400 578000
rect 475200 576000 475800 577400
rect 477200 576000 486400 577400
rect 475200 575400 486400 576000
rect 475200 574000 475800 575400
rect 477200 574000 486400 575400
rect 475200 573400 486400 574000
rect 475200 572000 475800 573400
rect 477200 572000 486400 573400
rect 475200 571400 486400 572000
rect 475200 570000 475800 571400
rect 477200 570400 486400 571400
rect 497000 584200 561400 594400
rect 497000 579200 503400 584200
rect 477200 570000 488400 570400
rect 475200 569400 488400 570000
rect 475200 568000 475800 569400
rect 477200 568000 488400 569400
rect 475200 567400 488400 568000
rect 475200 566000 475800 567400
rect 477200 566000 488400 567400
rect 475200 565400 488400 566000
rect 4400 562800 4800 564000
rect 6200 562800 7400 564000
rect 8800 562800 9200 564000
rect 4400 562000 9200 562800
rect 4400 560800 4800 562000
rect 6200 560800 7400 562000
rect 8800 560800 9200 562000
rect 4400 560000 9200 560800
rect 4400 558800 4800 560000
rect 6200 558800 7400 560000
rect 8800 558800 9200 560000
rect 4400 558000 9200 558800
rect 4400 556800 4800 558000
rect 6200 556800 7400 558000
rect 8800 556800 9200 558000
rect 4400 556000 9200 556800
rect 4400 554800 4800 556000
rect 6200 554800 7400 556000
rect 8800 554800 9200 556000
rect 4400 554000 9200 554800
rect 4400 552800 4800 554000
rect 6200 552800 7400 554000
rect 8800 552800 9200 554000
rect 4400 552000 9200 552800
rect 4400 550800 4800 552000
rect 6200 550800 7400 552000
rect 8800 550800 9200 552000
rect 4400 550000 9200 550800
rect 4400 548800 4800 550000
rect 6200 548800 7400 550000
rect 8800 548800 9200 550000
rect 4400 548000 9200 548800
rect 4400 546800 4800 548000
rect 6200 546800 7400 548000
rect 8800 546800 9200 548000
rect 4400 546000 9200 546800
rect 3200 544800 4800 546000
rect 6200 544800 7400 546000
rect 8800 544800 9200 546000
rect 3200 544000 9200 544800
rect 3200 542800 4800 544000
rect 6200 542800 7400 544000
rect 8800 542800 9200 544000
rect 3200 542000 9200 542800
rect 3200 540800 4800 542000
rect 6200 540800 7400 542000
rect 8800 540800 9200 542000
rect 3200 540000 9200 540800
rect 3200 538800 4800 540000
rect 6200 538800 7400 540000
rect 8800 538800 9200 540000
rect 3200 538000 9200 538800
rect 15400 564200 17400 564700
rect 15400 563600 16000 564200
rect 16800 563600 17400 564200
rect 15400 562200 15800 563600
rect 17000 562200 17400 563600
rect 15400 561600 17400 562200
rect 15400 560200 15800 561600
rect 17000 560200 17400 561600
rect 15400 559400 17400 560200
rect 15400 558000 15800 559400
rect 17000 558000 17400 559400
rect 15400 557600 16000 558000
rect 16800 557600 17400 558000
rect 15400 557200 17400 557600
rect 15400 555800 15800 557200
rect 17000 555800 17400 557200
rect 15400 555200 17400 555800
rect 15400 554800 16000 555200
rect 16800 554800 17400 555200
rect 15400 553400 15800 554800
rect 17000 553400 17400 554800
rect 15400 552600 17400 553400
rect 15400 551200 15800 552600
rect 17000 551200 17400 552600
rect 15400 550200 17400 551200
rect 15400 548800 15800 550200
rect 17000 548800 17400 550200
rect 15400 548600 16000 548800
rect 16800 548600 17400 548800
rect 15400 547800 17400 548600
rect 15400 547200 16000 547800
rect 16800 547200 17400 547800
rect 15400 544800 17400 547200
rect 15400 544200 16000 544800
rect 16800 544400 17400 544800
rect 475200 564000 475800 565400
rect 477200 564000 488400 565400
rect 475200 563400 488400 564000
rect 475200 562000 475800 563400
rect 477200 562000 488400 563400
rect 475200 561400 488400 562000
rect 475200 560000 475800 561400
rect 477200 560000 488400 561400
rect 475200 559400 488400 560000
rect 497000 567600 503200 579200
rect 549600 577400 561400 584200
rect 511690 574080 519090 574680
rect 504810 572500 505930 572580
rect 504810 572030 504870 572500
rect 505860 572030 505930 572500
rect 504810 571350 505930 572030
rect 504810 570440 504940 571350
rect 505850 570440 505930 571350
rect 504810 570360 505930 570440
rect 511690 568680 512590 574080
rect 518490 568680 519090 574080
rect 511690 567980 519090 568680
rect 529400 571400 539000 572400
rect 497000 564600 497200 567600
rect 502800 566600 503200 567600
rect 502800 564600 508000 566600
rect 497000 563000 508000 564600
rect 497000 560000 501400 563000
rect 507000 560000 508000 563000
rect 497000 559800 508000 560000
rect 475200 558000 475800 559400
rect 477200 558000 488400 559400
rect 475200 557400 488400 558000
rect 495460 557800 495700 557830
rect 475200 556000 475800 557400
rect 477200 556000 486400 557400
rect 495460 556610 495490 557800
rect 495680 557400 495700 557800
rect 500400 557400 508000 559800
rect 495680 557000 499790 557400
rect 495680 556610 495700 557000
rect 495460 556580 495700 556610
rect 475200 555400 486400 556000
rect 475200 554000 475800 555400
rect 477200 554000 486400 555400
rect 475200 553400 486400 554000
rect 475200 552000 475800 553400
rect 477200 552000 486400 553400
rect 475200 551400 486400 552000
rect 475200 550000 475800 551400
rect 477200 550000 486400 551400
rect 475200 549400 486400 550000
rect 475200 548000 475800 549400
rect 477200 548000 486400 549400
rect 475200 547400 486400 548000
rect 475200 546000 475800 547400
rect 477200 546000 486400 547400
rect 475200 545400 486400 546000
rect 475200 544400 475800 545400
rect 16800 544200 475800 544400
rect 15400 544000 475800 544200
rect 477200 544000 486400 545400
rect 15400 543400 486400 544000
rect 15400 542200 475800 543400
rect 15400 541800 17400 542200
rect 15400 541200 16000 541800
rect 16800 541200 17400 541800
rect 15400 538800 17400 541200
rect 15400 538200 16000 538800
rect 16800 538200 17400 538800
rect 3200 537600 5800 538000
rect 3200 536400 3800 537600
rect 5200 536590 5800 537600
rect 6880 536700 7340 536740
rect 6880 536590 6920 536700
rect 5200 536400 6920 536590
rect 3200 535600 6920 536400
rect 3200 534400 3800 535600
rect 5200 534760 6920 535600
rect 5200 534400 5800 534760
rect 6880 534720 6920 534760
rect 7200 534720 7340 536700
rect 6880 534680 7340 534720
rect 8380 536700 8740 536740
rect 8380 534720 8420 536700
rect 8700 536590 8740 536700
rect 15400 536590 17400 538200
rect 8700 535800 17400 536590
rect 8700 535200 16000 535800
rect 16800 535200 17400 535800
rect 8700 534790 17400 535200
rect 8700 534720 8740 534790
rect 8380 534680 8740 534720
rect 3200 533600 5800 534400
rect 3200 532400 3800 533600
rect 5200 532400 5800 533600
rect 10000 532800 10600 533200
rect 3200 532080 5800 532400
rect 3200 531700 3710 532080
rect 4140 531700 4930 532080
rect 5360 531700 5800 532080
rect 3200 531600 5800 531700
rect 3200 531120 3800 531600
rect 5200 531120 5800 531600
rect 3200 530740 3700 531120
rect 5350 530740 5800 531120
rect 3200 530400 3800 530740
rect 5200 530400 5800 530740
rect 3200 530170 5800 530400
rect 3200 529790 3660 530170
rect 4090 529790 4880 530170
rect 5310 529790 5800 530170
rect 3200 529600 5800 529790
rect 3200 529050 3800 529600
rect 5200 529050 5800 529600
rect 3200 528670 3700 529050
rect 5350 528670 5800 529050
rect 3200 528400 3800 528670
rect 5200 528400 5800 528670
rect 3200 528180 5800 528400
rect 3200 527800 3680 528180
rect 4110 527800 4900 528180
rect 5330 527800 5800 528180
rect 3200 527600 5800 527800
rect 3200 526400 3800 527600
rect 5200 526400 5800 527600
rect 15400 532200 17400 534790
rect 15400 531800 15800 532200
rect 17100 531800 17400 532200
rect 15400 531500 17400 531800
rect 15400 531100 15800 531500
rect 17100 531100 17400 531500
rect 15400 530900 17400 531100
rect 15400 530500 15800 530900
rect 17100 530500 17400 530900
rect 15400 530200 17400 530500
rect 15400 529800 15800 530200
rect 17100 529800 17400 530200
rect 15400 529500 17400 529800
rect 15400 529100 15800 529500
rect 17100 529100 17400 529500
rect 15400 528800 17400 529100
rect 15400 528400 15800 528800
rect 17100 528400 17400 528800
rect 10000 527000 10600 527400
rect 15400 527200 17400 528400
rect 3200 525600 5800 526400
rect 3200 524400 3800 525600
rect 5200 524400 5800 525600
rect 3200 523600 5800 524400
rect 3200 522400 3800 523600
rect 5200 522400 5800 523600
rect 3200 521600 5800 522400
rect 3200 520400 3800 521600
rect 5200 520400 5800 521600
rect 3200 519600 5800 520400
rect 3200 518400 3800 519600
rect 5200 518400 5800 519600
rect 3200 517600 5800 518400
rect 3200 516400 3800 517600
rect 5200 516400 5800 517600
rect 3200 515600 5800 516400
rect 3200 514400 3800 515600
rect 5200 514400 5800 515600
rect 3200 513600 5800 514400
rect 3200 512400 3800 513600
rect 5200 512400 5800 513600
rect 3200 511600 5800 512400
rect 3200 510400 3800 511600
rect 5200 510400 5800 511600
rect 3200 509600 5800 510400
rect 3200 508400 3800 509600
rect 5200 508400 5800 509600
rect 3200 507600 5800 508400
rect 3200 506400 3800 507600
rect 5200 506400 5800 507600
rect 3200 505600 5800 506400
rect 3200 504400 3800 505600
rect 5200 504400 5800 505600
rect 3200 503600 5800 504400
rect 3200 502400 3800 503600
rect 5200 502400 5800 503600
rect 3200 501600 5800 502400
rect 3200 500400 3800 501600
rect 5200 500400 5800 501600
rect 3200 499600 5800 500400
rect 3200 498400 3800 499600
rect 5200 498400 5800 499600
rect 3200 497600 5800 498400
rect 3200 496400 3800 497600
rect 5200 496400 5800 497600
rect 3200 495600 5800 496400
rect 3200 494400 3800 495600
rect 5200 494400 5800 495600
rect 3200 493600 5800 494400
rect 3200 492400 3800 493600
rect 5200 492400 5800 493600
rect 3200 491600 5800 492400
rect 3200 490400 3800 491600
rect 5200 490400 5800 491600
rect 3200 489600 5800 490400
rect 3200 488400 3800 489600
rect 5200 488400 5800 489600
rect 3200 487600 5800 488400
rect 3200 486400 3800 487600
rect 5200 486400 5800 487600
rect 3200 485600 5800 486400
rect 3200 484400 3800 485600
rect 5200 484400 5800 485600
rect 3200 483600 5800 484400
rect 3200 482400 3800 483600
rect 5200 482400 5800 483600
rect 3200 481600 5800 482400
rect 3200 480400 3800 481600
rect 5200 480400 5800 481600
rect 3200 479600 5800 480400
rect 3200 478400 3800 479600
rect 5200 478400 5800 479600
rect 3200 477600 5800 478400
rect 3200 476400 3800 477600
rect 5200 476400 5800 477600
rect 3200 475600 5800 476400
rect 3200 474400 3800 475600
rect 5200 474400 5800 475600
rect 3200 473600 5800 474400
rect 3200 472400 3800 473600
rect 5200 472400 5800 473600
rect 3200 471600 5800 472400
rect 3200 470400 3800 471600
rect 5200 470400 5800 471600
rect 3200 469600 5800 470400
rect 3200 468400 3800 469600
rect 5200 468400 5800 469600
rect 3200 467600 5800 468400
rect 3200 466400 3800 467600
rect 5200 466400 5800 467600
rect 3200 465600 5800 466400
rect 3200 464400 3800 465600
rect 5200 464400 5800 465600
rect 3200 463600 5800 464400
rect 3200 462400 3800 463600
rect 5200 462400 5800 463600
rect 3200 461600 5800 462400
rect 3200 460400 3800 461600
rect 5200 460400 5800 461600
rect 3200 459600 5800 460400
rect 3200 458400 3800 459600
rect 5200 458400 5800 459600
rect 3200 457600 5800 458400
rect 3200 456400 3800 457600
rect 5200 456400 5800 457600
rect 3200 455600 5800 456400
rect 3200 454400 3800 455600
rect 5200 454400 5800 455600
rect 3200 453600 5800 454400
rect 3200 452400 3800 453600
rect 5200 452400 5800 453600
rect 3200 451600 5800 452400
rect 3200 450400 3800 451600
rect 5200 450400 5800 451600
rect 3200 449600 5800 450400
rect 3200 448400 3800 449600
rect 5200 448400 5800 449600
rect 3200 447600 5800 448400
rect 3200 446400 3800 447600
rect 5200 446400 5800 447600
rect 3200 445600 5800 446400
rect 3200 444400 3800 445600
rect 5200 444400 5800 445600
rect 3200 443600 5800 444400
rect 3200 442400 3800 443600
rect 5200 442400 5800 443600
rect 3200 441600 5800 442400
rect 3200 440400 3800 441600
rect 5200 440400 5800 441600
rect 3200 439600 5800 440400
rect 3200 438400 3800 439600
rect 5200 438400 5800 439600
rect 3200 437600 5800 438400
rect 3200 436400 3800 437600
rect 5200 436400 5800 437600
rect 3200 435600 5800 436400
rect 3200 434400 3800 435600
rect 5200 434400 5800 435600
rect 3200 433600 5800 434400
rect 3200 432400 3800 433600
rect 5200 432400 5800 433600
rect 3200 431000 5800 432400
rect 15400 526600 16000 527200
rect 16800 526600 17400 527200
rect 15400 524200 17400 526600
rect 15400 523600 16000 524200
rect 16800 523600 17400 524200
rect 15400 521200 17400 523600
rect 15400 520600 16000 521200
rect 16800 520600 17400 521200
rect 15400 518200 17400 520600
rect 15400 517600 16000 518200
rect 16800 517600 17400 518200
rect 15400 515200 17400 517600
rect 15400 514600 16000 515200
rect 16800 514600 17400 515200
rect 15400 512200 17400 514600
rect 15400 511600 16000 512200
rect 16800 511600 17400 512200
rect 15400 509200 17400 511600
rect 15400 508600 16000 509200
rect 16800 508600 17400 509200
rect 15400 506200 17400 508600
rect 15400 505600 16000 506200
rect 16800 505600 17400 506200
rect 15400 503200 17400 505600
rect 15400 502600 16000 503200
rect 16800 502600 17400 503200
rect 15400 500200 17400 502600
rect 15400 499600 16000 500200
rect 16800 499600 17400 500200
rect 15400 497200 17400 499600
rect 15400 496600 16000 497200
rect 16800 496600 17400 497200
rect 15400 494200 17400 496600
rect 15400 493600 16000 494200
rect 16800 493600 17400 494200
rect 15400 491200 17400 493600
rect 15400 490600 16000 491200
rect 16800 490600 17400 491200
rect 15400 488200 17400 490600
rect 15400 487600 16000 488200
rect 16800 487600 17400 488200
rect 15400 485200 17400 487600
rect 15400 484600 16000 485200
rect 16800 484600 17400 485200
rect 15400 482200 17400 484600
rect 15400 481600 16000 482200
rect 16800 481600 17400 482200
rect 15400 479200 17400 481600
rect 15400 478600 16000 479200
rect 16800 478600 17400 479200
rect 15400 476200 17400 478600
rect 15400 475600 16000 476200
rect 16800 475600 17400 476200
rect 15400 473200 17400 475600
rect 15400 472600 16000 473200
rect 16800 472600 17400 473200
rect 15400 470200 17400 472600
rect 15400 469600 16000 470200
rect 16800 469600 17400 470200
rect 15400 467200 17400 469600
rect 15400 466600 16000 467200
rect 16800 466600 17400 467200
rect 15400 464200 17400 466600
rect 15400 463600 16000 464200
rect 16800 463600 17400 464200
rect 15400 461200 17400 463600
rect 15400 460600 16000 461200
rect 16800 460600 17400 461200
rect 15400 458200 17400 460600
rect 15400 457600 16000 458200
rect 16800 457600 17400 458200
rect 15400 455200 17400 457600
rect 15400 454600 16000 455200
rect 16800 454600 17400 455200
rect 15400 452200 17400 454600
rect 15400 451600 16000 452200
rect 16800 451600 17400 452200
rect 15400 449200 17400 451600
rect 15400 448600 16000 449200
rect 16800 448600 17400 449200
rect 15400 446200 17400 448600
rect 15400 445600 16000 446200
rect 16800 445600 17400 446200
rect 15400 443200 17400 445600
rect 15400 442600 16000 443200
rect 16800 442600 17400 443200
rect 15400 440200 17400 442600
rect 15400 439600 16000 440200
rect 16800 439600 17400 440200
rect 15400 437200 17400 439600
rect 15400 436600 16000 437200
rect 16800 436600 17400 437200
rect 15400 434200 17400 436600
rect 15400 433600 16000 434200
rect 16800 433600 17400 434200
rect 15400 431200 17400 433600
rect 15400 430600 16000 431200
rect 16800 430600 17400 431200
rect 15400 428200 17400 430600
rect 15400 427600 16000 428200
rect 16800 427600 17400 428200
rect 15400 425200 17400 427600
rect 15400 424600 16000 425200
rect 16800 424600 17400 425200
rect 15400 422200 17400 424600
rect 15400 421600 16000 422200
rect 16800 421600 17400 422200
rect 15400 419200 17400 421600
rect 15400 418600 16000 419200
rect 16800 418600 17400 419200
rect 15400 416200 17400 418600
rect 15400 415600 16000 416200
rect 16800 415600 17400 416200
rect 15400 413200 17400 415600
rect 15400 412600 16000 413200
rect 16800 412600 17400 413200
rect 15400 410200 17400 412600
rect 15400 409600 16000 410200
rect 16800 409600 17400 410200
rect 15400 407200 17400 409600
rect 15400 406600 16000 407200
rect 16800 406600 17400 407200
rect 15400 404200 17400 406600
rect 15400 403600 16000 404200
rect 16800 403600 17400 404200
rect 15400 401200 17400 403600
rect 15400 400600 16000 401200
rect 16800 400600 17400 401200
rect 15400 398200 17400 400600
rect 15400 397600 16000 398200
rect 16800 397600 17400 398200
rect 15400 395200 17400 397600
rect 15400 394600 16000 395200
rect 16800 394600 17400 395200
rect 15400 392200 17400 394600
rect 15400 391600 16000 392200
rect 16800 391600 17400 392200
rect 15400 389200 17400 391600
rect 15400 388600 16000 389200
rect 16800 388600 17400 389200
rect 15400 386200 17400 388600
rect 15400 385600 16000 386200
rect 16800 385600 17400 386200
rect 15400 383200 17400 385600
rect 15400 382600 16000 383200
rect 16800 382600 17400 383200
rect 15400 380200 17400 382600
rect 15400 379600 16000 380200
rect 16800 379600 17400 380200
rect 15400 377200 17400 379600
rect 15400 376600 16000 377200
rect 16800 376600 17400 377200
rect 600 375400 2400 375600
rect 600 375000 1000 375400
rect 2000 375000 2400 375400
rect 600 374800 2400 375000
rect 600 374400 1000 374800
rect 2000 374400 2400 374800
rect 600 374000 2400 374400
rect 600 373600 1000 374000
rect 2000 373600 2400 374000
rect 600 373200 2400 373600
rect 600 372800 1000 373200
rect 2000 372800 2400 373200
rect 600 372400 2400 372800
rect 600 372000 1000 372400
rect 2000 372000 2400 372400
rect 600 371600 2400 372000
rect 600 371200 1000 371600
rect 2000 371200 2400 371600
rect 600 370800 2400 371200
rect 600 370400 1000 370800
rect 2000 370400 2400 370800
rect 600 370000 2400 370400
rect 15400 374200 17400 376600
rect 15400 373600 16000 374200
rect 16800 373600 17400 374200
rect 15400 371200 17400 373600
rect 15400 370600 16000 371200
rect 16800 370600 17400 371200
rect 600 369400 1600 370000
rect 600 368800 800 369400
rect 1400 368800 1600 369400
rect 600 367400 1600 368800
rect 600 366800 800 367400
rect 1400 366800 1600 367400
rect 2000 368190 3100 368200
rect 2000 368000 10573 368190
rect 2000 367200 2700 368000
rect 10400 367200 10573 368000
rect 2000 367070 10573 367200
rect 15400 367100 17400 370600
rect 2000 367000 6583 367070
rect 600 365400 1600 366800
rect 600 364800 800 365400
rect 1400 364800 1600 365400
rect 600 363400 1600 364800
rect 600 362800 800 363400
rect 1400 362800 1600 363400
rect 600 361400 1600 362800
rect 600 360800 800 361400
rect 1400 360800 1600 361400
rect 600 359400 1600 360800
rect 600 358800 800 359400
rect 1400 358800 1600 359400
rect 600 357400 1600 358800
rect 600 356800 800 357400
rect 1400 356800 1600 357400
rect 600 355400 1600 356800
rect 600 354800 800 355400
rect 1400 354800 1600 355400
rect 600 353400 1600 354800
rect 600 352800 800 353400
rect 1400 352800 1600 353400
rect 600 351400 1600 352800
rect 600 350800 800 351400
rect 1400 350800 1600 351400
rect 600 349400 1600 350800
rect 600 348800 800 349400
rect 1400 348800 1600 349400
rect 600 347400 1600 348800
rect 600 346800 800 347400
rect 1400 346800 1600 347400
rect 600 345400 1600 346800
rect 600 344800 800 345400
rect 1400 344800 1600 345400
rect 600 344200 1600 344800
rect 2013 366990 6583 367000
rect 2013 344290 2133 366990
rect 15400 366800 15800 367100
rect 17100 366800 17400 367100
rect 15400 366100 17400 366800
rect 15400 365800 15800 366100
rect 17100 365800 17400 366100
rect 15400 365100 17400 365800
rect 15400 364800 15800 365100
rect 17100 364800 17400 365100
rect 15400 364100 17400 364800
rect 15400 363800 15800 364100
rect 17100 363800 17400 364100
rect 15400 363100 17400 363800
rect 15400 362800 15800 363100
rect 17100 362800 17400 363100
rect 15400 362100 17400 362800
rect 15400 361800 15800 362100
rect 17100 361800 17400 362100
rect 15400 361100 17400 361800
rect 15400 360800 15800 361100
rect 17100 360800 17400 361100
rect 15400 360100 17400 360800
rect 15400 359800 15800 360100
rect 17100 359800 17400 360100
rect 15400 359100 17400 359800
rect 15400 358800 15800 359100
rect 17100 358800 17400 359100
rect 15400 358100 17400 358800
rect 15400 357800 15800 358100
rect 17100 357800 17400 358100
rect 15400 357100 17400 357800
rect 15400 356800 15800 357100
rect 17100 356800 17400 357100
rect 15400 356100 17400 356800
rect 15400 355800 15800 356100
rect 17100 355800 17400 356100
rect 15400 355100 17400 355800
rect 15400 354800 15800 355100
rect 17100 354800 17400 355100
rect 15400 354100 17400 354800
rect 15400 353800 15800 354100
rect 17100 353800 17400 354100
rect 15400 353100 17400 353800
rect 15400 352800 15800 353100
rect 17100 352800 17400 353100
rect 15400 352100 17400 352800
rect 15400 351800 15800 352100
rect 17100 351800 17400 352100
rect 15400 351100 17400 351800
rect 15400 350800 15800 351100
rect 17100 350800 17400 351100
rect 15400 350100 17400 350800
rect 15400 349800 15800 350100
rect 17100 349800 17400 350100
rect 15400 349100 17400 349800
rect 15400 348800 15800 349100
rect 17100 348800 17400 349100
rect 15400 348100 17400 348800
rect 15400 347800 15800 348100
rect 17100 347800 17400 348100
rect 15400 347100 17400 347800
rect 15400 346800 15800 347100
rect 17100 346800 17400 347100
rect 15400 346100 17400 346800
rect 15400 345800 15800 346100
rect 17100 345800 17400 346100
rect 15400 345100 17400 345800
rect 15400 344800 15800 345100
rect 17100 344800 17400 345100
rect 6103 344680 6343 344710
rect 6103 344290 6123 344680
rect 2013 343890 6123 344290
rect 6103 343490 6123 343890
rect 6313 343490 6343 344680
rect 6103 343460 6343 343490
rect 15400 344100 17400 344800
rect 15400 343800 15800 344100
rect 17100 343800 17400 344100
rect 15400 341800 17400 343800
rect 15400 341200 16000 341800
rect 16800 341200 17400 341800
rect 15400 341100 17400 341200
rect 12900 340600 17400 341100
rect 12900 340300 13800 340600
rect 15000 340300 17400 340600
rect 12900 339600 17400 340300
rect 12900 339300 13800 339600
rect 15000 339300 17400 339600
rect 12900 338800 17400 339300
rect 12900 338600 16000 338800
rect 12900 338300 13800 338600
rect 15000 338300 16000 338600
rect 12900 338200 16000 338300
rect 16800 338200 17400 338800
rect 12900 337600 17400 338200
rect 12900 337300 13800 337600
rect 15000 337300 17400 337600
rect 12900 336600 17400 337300
rect 12900 336300 13800 336600
rect 15000 336300 17400 336600
rect 12900 335800 17400 336300
rect 12900 335600 16000 335800
rect 12900 335300 13800 335600
rect 15000 335300 16000 335600
rect 12900 335200 16000 335300
rect 16800 335200 17400 335800
rect 12900 334600 17400 335200
rect 12900 334300 13800 334600
rect 15000 334300 17400 334600
rect 12900 333600 17400 334300
rect 12900 333300 13800 333600
rect 15000 333300 17400 333600
rect 12900 333000 17400 333300
rect 15400 332800 17400 333000
rect 15400 332200 16000 332800
rect 16800 332200 17400 332800
rect 15400 331400 17400 332200
rect 475200 542000 475800 542200
rect 477200 542000 486400 543400
rect 475200 541400 486400 542000
rect 475200 540000 475800 541400
rect 477200 540000 486400 541400
rect 475200 539400 486400 540000
rect 475200 538000 475800 539400
rect 477200 538000 486400 539400
rect 475200 537400 486400 538000
rect 475200 536000 475800 537400
rect 477200 536000 486400 537400
rect 475200 535400 486400 536000
rect 475200 534000 475800 535400
rect 477200 534000 486400 535400
rect 499670 534300 499790 557000
rect 500400 554400 501400 557400
rect 507000 554400 508000 557400
rect 500400 550000 508000 554400
rect 529400 558400 541000 571400
rect 549600 567600 555800 577400
rect 564280 574210 571680 574810
rect 557400 572630 558520 572710
rect 557400 572160 557460 572630
rect 558450 572160 558520 572630
rect 557400 571230 558520 572160
rect 557400 570740 557670 571230
rect 558130 570740 558520 571230
rect 557400 570600 558520 570740
rect 564280 568810 565180 574210
rect 571080 568810 571680 574210
rect 564280 568110 571680 568810
rect 549600 564600 549800 567600
rect 555400 566800 555800 567600
rect 555400 564600 560400 566800
rect 549600 563600 560400 564600
rect 549600 560600 553800 563600
rect 559400 560600 560400 563600
rect 549600 560000 560400 560600
rect 529400 554200 539000 558400
rect 552800 558000 560400 560000
rect 548050 557930 548290 557960
rect 548050 556740 548080 557930
rect 548270 557530 548290 557930
rect 548270 557130 552380 557530
rect 548270 556740 548290 557130
rect 548050 556710 548290 556740
rect 500400 547000 501400 550000
rect 507000 547000 508000 550000
rect 500400 544200 508000 547000
rect 511790 551080 519190 551780
rect 511790 545680 512790 551080
rect 518690 545680 519190 551080
rect 511790 545080 519190 545680
rect 500400 541200 501400 544200
rect 507000 541200 508000 544200
rect 500400 538400 508000 541200
rect 500400 535400 501400 538400
rect 507000 535400 508000 538400
rect 500400 534800 508000 535400
rect 495220 534220 499790 534300
rect 475200 533800 486400 534000
rect 491230 533910 499790 534220
rect 491230 533850 499110 533910
rect 475200 533400 485800 533800
rect 475200 532000 475800 533400
rect 477200 532000 485800 533400
rect 475200 531400 485800 532000
rect 491230 532700 491350 533850
rect 499020 532700 499110 533850
rect 491230 531460 499110 532700
rect 527800 533600 539000 554200
rect 552260 534430 552380 557130
rect 552800 555000 553800 558000
rect 559400 555000 560400 558000
rect 552800 550600 560400 555000
rect 552800 547600 553800 550600
rect 559400 547600 560400 550600
rect 552800 544800 560400 547600
rect 564380 551210 571780 551910
rect 564380 545810 565380 551210
rect 571280 545810 571780 551210
rect 564380 545210 571780 545810
rect 552800 541800 553800 544800
rect 559400 541800 560400 544800
rect 552800 540200 560400 541800
rect 575600 540200 582600 540400
rect 552800 539000 582600 540200
rect 552800 536000 553800 539000
rect 559400 536000 582600 539000
rect 552800 535200 582600 536000
rect 547810 534350 552380 534430
rect 543820 534040 552380 534350
rect 543820 533980 551700 534040
rect 475200 530000 475800 531400
rect 477200 530000 485800 531400
rect 475200 529400 485800 530000
rect 475200 528000 475800 529400
rect 477200 528000 485800 529400
rect 475200 527400 485800 528000
rect 475200 526000 475800 527400
rect 477200 526000 485800 527400
rect 475200 525400 485800 526000
rect 475200 524000 475800 525400
rect 477200 524000 485800 525400
rect 475200 523400 485800 524000
rect 475200 522000 475800 523400
rect 477200 522000 485800 523400
rect 475200 521400 485800 522000
rect 475200 520000 475800 521400
rect 477200 520000 485800 521400
rect 511890 527380 519190 528080
rect 511890 522080 512590 527380
rect 518590 522080 519190 527380
rect 511890 521380 519190 522080
rect 475200 519400 485800 520000
rect 475200 518000 475800 519400
rect 477200 518000 485800 519400
rect 475200 517400 485800 518000
rect 475200 516000 475800 517400
rect 477200 516200 485800 517400
rect 527800 516200 537400 533600
rect 543820 532830 543940 533980
rect 551610 532830 551700 533980
rect 557800 533200 582600 535200
rect 543820 531590 551700 532830
rect 564480 527510 571780 528210
rect 564480 522210 565180 527510
rect 571180 522210 571780 527510
rect 564480 521510 571780 522210
rect 477200 516000 537400 516200
rect 475200 515400 537400 516000
rect 475200 514000 475800 515400
rect 477200 514000 567600 515400
rect 575600 515200 582600 533200
rect 475200 513400 567600 514000
rect 475200 512000 475800 513400
rect 477200 512000 567600 513400
rect 475200 511400 567600 512000
rect 475200 510000 475800 511400
rect 477200 510000 567600 511400
rect 475200 509400 567600 510000
rect 475200 508000 475800 509400
rect 477200 508000 567600 509400
rect 475200 507400 567600 508000
rect 475200 506000 475800 507400
rect 477200 506600 567600 507400
rect 477200 506000 477800 506600
rect 475200 505400 477800 506000
rect 530400 505800 567600 506600
rect 475200 504000 475800 505400
rect 477200 504000 477800 505400
rect 475200 503400 477800 504000
rect 554600 503800 567600 505800
rect 571200 504800 582600 515200
rect 475200 502000 475800 503400
rect 477200 502000 477800 503400
rect 475200 501400 477800 502000
rect 475200 500000 475800 501400
rect 477200 500000 477800 501400
rect 475200 499400 477800 500000
rect 475200 498000 475800 499400
rect 477200 498000 477800 499400
rect 475200 497400 477800 498000
rect 475200 496000 475800 497400
rect 477200 496000 477800 497400
rect 475200 495400 477800 496000
rect 475200 494000 475800 495400
rect 477200 494000 477800 495400
rect 475200 493400 477800 494000
rect 475200 492000 475800 493400
rect 477200 492000 477800 493400
rect 528170 500750 530930 500870
rect 528170 493080 529410 500750
rect 530560 496880 530930 500750
rect 530560 493080 531010 496880
rect 553290 496610 554540 496640
rect 553290 496420 553320 496610
rect 554510 496420 554540 496610
rect 553290 496400 554540 496420
rect 528170 492990 531010 493080
rect 530620 492430 531010 492990
rect 553710 492430 554110 496400
rect 571200 494600 579400 504800
rect 530620 492310 554110 492430
rect 556800 494400 579400 494600
rect 556800 494200 562000 494400
rect 475200 491400 477800 492000
rect 556800 491600 557800 494200
rect 475200 490000 475800 491400
rect 477200 490000 477800 491400
rect 475200 489400 477800 490000
rect 475200 488000 475800 489400
rect 477200 488000 477800 489400
rect 475200 487400 477800 488000
rect 475200 486000 475800 487400
rect 477200 486000 477800 487400
rect 475200 485400 477800 486000
rect 475200 484000 475800 485400
rect 477200 484000 477800 485400
rect 528400 490600 557800 491600
rect 528400 485000 529000 490600
rect 532000 485000 534800 490600
rect 537800 485000 540600 490600
rect 543600 485000 548000 490600
rect 551000 485000 553600 490600
rect 556600 488600 557800 490600
rect 560800 488800 562000 494200
rect 565000 488800 579400 494400
rect 560800 488600 579400 488800
rect 556600 488000 571000 488600
rect 556600 485000 559800 488000
rect 567070 487230 569290 487290
rect 567070 487160 568740 487230
rect 567070 486250 567150 487160
rect 568060 486250 568740 487160
rect 567070 486240 568740 486250
rect 569210 486240 569290 487230
rect 567070 486170 569290 486240
rect 528400 484000 559800 485000
rect 475200 483400 477800 484000
rect 475200 482000 475800 483400
rect 477200 482000 477800 483400
rect 475200 481400 477800 482000
rect 475200 480000 475800 481400
rect 477200 480000 477800 481400
rect 475200 479400 477800 480000
rect 475200 478000 475800 479400
rect 477200 478000 477800 479400
rect 475200 477400 477800 478000
rect 475200 476000 475800 477400
rect 477200 476000 477800 477400
rect 475200 475400 477800 476000
rect 475200 474000 475800 475400
rect 477200 474000 477800 475400
rect 475200 473400 477800 474000
rect 475200 472000 475800 473400
rect 477200 472000 477800 473400
rect 518090 479510 524790 480210
rect 518090 473510 518790 479510
rect 524090 473510 524790 479510
rect 518090 472910 524790 473510
rect 541790 479310 548490 480310
rect 541790 473410 542390 479310
rect 547790 473410 548490 479310
rect 541790 472910 548490 473410
rect 564690 479510 571390 480410
rect 564690 473610 565390 479510
rect 570790 473610 571390 479510
rect 564690 473010 571390 473610
rect 475200 471400 477800 472000
rect 475200 470000 475800 471400
rect 477200 470000 477800 471400
rect 475200 469400 477800 470000
rect 475200 468000 475800 469400
rect 477200 468000 477800 469400
rect 576200 468600 579400 488600
rect 475200 467400 477800 468000
rect 475200 466000 475800 467400
rect 477200 466000 477800 467400
rect 475200 465400 477800 466000
rect 475200 464000 475800 465400
rect 477200 464000 477800 465400
rect 475200 463400 477800 464000
rect 475200 462000 475800 463400
rect 477200 462000 477800 463400
rect 475200 461400 477800 462000
rect 475200 460000 475800 461400
rect 477200 460000 477800 461400
rect 475200 459400 477800 460000
rect 475200 458000 475800 459400
rect 477200 458000 477800 459400
rect 475200 457400 477800 458000
rect 475200 456000 475800 457400
rect 477200 456000 477800 457400
rect 475200 455400 477800 456000
rect 475200 454000 475800 455400
rect 477200 454000 477800 455400
rect 475200 453400 477800 454000
rect 475200 452000 475800 453400
rect 477200 452000 477800 453400
rect 475200 451400 477800 452000
rect 475200 450000 475800 451400
rect 477200 450000 477800 451400
rect 475200 449400 477800 450000
rect 475200 448000 475800 449400
rect 477200 448000 477800 449400
rect 475200 447400 477800 448000
rect 475200 446000 475800 447400
rect 477200 446000 477800 447400
rect 475200 445400 477800 446000
rect 475200 444000 475800 445400
rect 477200 444000 477800 445400
rect 475200 443400 477800 444000
rect 475200 442000 475800 443400
rect 477200 442000 477800 443400
rect 475200 441400 477800 442000
rect 475200 440000 475800 441400
rect 477200 440000 477800 441400
rect 475200 439400 477800 440000
rect 475200 438000 475800 439400
rect 477200 438000 477800 439400
rect 475200 437400 477800 438000
rect 475200 436000 475800 437400
rect 477200 436000 477800 437400
rect 475200 435400 477800 436000
rect 475200 434000 475800 435400
rect 477200 434000 477800 435400
rect 475200 433400 477800 434000
rect 475200 432000 475800 433400
rect 477200 432000 477800 433400
rect 475200 431400 477800 432000
rect 475200 430000 475800 431400
rect 477200 430000 477800 431400
rect 475200 429400 477800 430000
rect 475200 428000 475800 429400
rect 477200 428000 477800 429400
rect 475200 427400 477800 428000
rect 475200 426000 475800 427400
rect 477200 426000 477800 427400
rect 475200 425400 477800 426000
rect 475200 424000 475800 425400
rect 477200 424000 477800 425400
rect 475200 423400 477800 424000
rect 475200 422000 475800 423400
rect 477200 422000 477800 423400
rect 475200 421400 477800 422000
rect 475200 420000 475800 421400
rect 477200 420000 477800 421400
rect 475200 419400 477800 420000
rect 475200 418000 475800 419400
rect 477200 418000 477800 419400
rect 475200 417400 477800 418000
rect 475200 416000 475800 417400
rect 477200 416000 477800 417400
rect 475200 415400 477800 416000
rect 475200 414000 475800 415400
rect 477200 414000 477800 415400
rect 475200 413400 477800 414000
rect 475200 412000 475800 413400
rect 477200 412000 477800 413400
rect 475200 411400 477800 412000
rect 475200 410000 475800 411400
rect 477200 410000 477800 411400
rect 475200 409400 477800 410000
rect 475200 408000 475800 409400
rect 477200 408000 477800 409400
rect 475200 407400 477800 408000
rect 475200 406000 475800 407400
rect 477200 406000 477800 407400
rect 475200 405400 477800 406000
rect 475200 404000 475800 405400
rect 477200 404000 477800 405400
rect 475200 403400 477800 404000
rect 475200 402000 475800 403400
rect 477200 402000 477800 403400
rect 475200 401400 477800 402000
rect 475200 400000 475800 401400
rect 477200 400000 477800 401400
rect 475200 399400 477800 400000
rect 475200 398000 475800 399400
rect 477200 398000 477800 399400
rect 475200 397400 477800 398000
rect 475200 396000 475800 397400
rect 477200 396000 477800 397400
rect 475200 395400 477800 396000
rect 475200 394000 475800 395400
rect 477200 394000 477800 395400
rect 475200 393400 477800 394000
rect 475200 392000 475800 393400
rect 477200 392000 477800 393400
rect 475200 391400 477800 392000
rect 475200 390000 475800 391400
rect 477200 390000 477800 391400
rect 475200 389400 477800 390000
rect 475200 388000 475800 389400
rect 477200 388000 477800 389400
rect 475200 387400 477800 388000
rect 475200 386000 475800 387400
rect 477200 386000 477800 387400
rect 475200 385400 477800 386000
rect 475200 384000 475800 385400
rect 477200 384000 477800 385400
rect 475200 383400 477800 384000
rect 475200 382000 475800 383400
rect 477200 382000 477800 383400
rect 475200 381400 477800 382000
rect 475200 380000 475800 381400
rect 477200 380000 477800 381400
rect 475200 379400 477800 380000
rect 475200 378000 475800 379400
rect 477200 378000 477800 379400
rect 475200 377400 477800 378000
rect 475200 376000 475800 377400
rect 477200 376000 477800 377400
rect 475200 375400 477800 376000
rect 475200 374000 475800 375400
rect 477200 374000 477800 375400
rect 475200 373400 477800 374000
rect 475200 372000 475800 373400
rect 477200 372000 477800 373400
rect 475200 371400 477800 372000
rect 475200 370000 475800 371400
rect 477200 370000 477800 371400
rect 475200 369400 477800 370000
rect 475200 368000 475800 369400
rect 477200 368000 477800 369400
rect 475200 367400 477800 368000
rect 475200 366000 475800 367400
rect 477200 366000 477800 367400
rect 475200 365400 477800 366000
rect 475200 364000 475800 365400
rect 477200 364000 477800 365400
rect 475200 363400 477800 364000
rect 475200 362000 475800 363400
rect 477200 362000 477800 363400
rect 475200 361400 477800 362000
rect 475200 360000 475800 361400
rect 477200 360000 477800 361400
rect 475200 359400 477800 360000
rect 475200 358000 475800 359400
rect 477200 358000 477800 359400
rect 475200 357400 477800 358000
rect 475200 356000 475800 357400
rect 477200 356000 477800 357400
rect 475200 355400 477800 356000
rect 475200 354000 475800 355400
rect 477200 354000 477800 355400
rect 475200 353400 477800 354000
rect 475200 352000 475800 353400
rect 477200 352000 477800 353400
rect 475200 351400 477800 352000
rect 475200 350000 475800 351400
rect 477200 350000 477800 351400
rect 475200 349400 477800 350000
rect 475200 348000 475800 349400
rect 477200 348000 477800 349400
rect 475200 347400 477800 348000
rect 475200 346000 475800 347400
rect 477200 346000 477800 347400
rect 475200 345400 477800 346000
rect 475200 344000 475800 345400
rect 477200 344000 477800 345400
rect 475200 343400 477800 344000
rect 475200 342000 475800 343400
rect 477200 342000 477800 343400
rect 475200 341400 477800 342000
rect 475200 340000 475800 341400
rect 477200 340000 477800 341400
rect 475200 339400 477800 340000
rect 475200 338000 475800 339400
rect 477200 338000 477800 339400
rect 475200 337400 477800 338000
rect 475200 336000 475800 337400
rect 477200 336000 477800 337400
rect 475200 335400 477800 336000
rect 475200 334000 475800 335400
rect 477200 334000 477800 335400
rect 475200 333400 477800 334000
rect 475200 332000 475800 333400
rect 477200 332000 477800 333400
rect 475200 331400 477800 332000
rect 15800 329800 17000 331400
rect 15800 329200 16000 329800
rect 16800 329200 17000 329800
rect 15800 326800 17000 329200
rect 4150 326173 6260 326233
rect 4150 325963 5710 326173
rect 4150 325503 4290 325963
rect 4780 325503 5710 325963
rect 4150 325183 5710 325503
rect 6180 325183 6260 326173
rect 4150 325113 6260 325183
rect 15800 326200 16000 326800
rect 16800 326200 17000 326800
rect 15800 323800 17000 326200
rect 15800 323200 16000 323800
rect 16800 323200 17000 323800
rect 15800 320800 17000 323200
rect 15800 320200 16000 320800
rect 16800 320200 17000 320800
rect 15800 317800 17000 320200
rect 15800 317200 16000 317800
rect 16800 317200 17000 317800
rect 15800 314800 17000 317200
rect 15800 314200 16000 314800
rect 16800 314200 17000 314800
rect 15800 311800 17000 314200
rect 15800 311200 16000 311800
rect 16800 311200 17000 311800
rect 15800 308800 17000 311200
rect 15800 308200 16000 308800
rect 16800 308200 17000 308800
rect 15800 305800 17000 308200
rect 15800 305200 16000 305800
rect 16800 305200 17000 305800
rect 15800 302800 17000 305200
rect 15800 302200 16000 302800
rect 16800 302200 17000 302800
rect 15800 299800 17000 302200
rect 15800 299200 16000 299800
rect 16800 299200 17000 299800
rect 15800 296800 17000 299200
rect 15800 296200 16000 296800
rect 16800 296200 17000 296800
rect 15800 293800 17000 296200
rect 15800 293200 16000 293800
rect 16800 293200 17000 293800
rect 15800 290800 17000 293200
rect 15800 290200 16000 290800
rect 16800 290200 17000 290800
rect 15800 287800 17000 290200
rect 15800 287200 16000 287800
rect 16800 287200 17000 287800
rect 15800 284800 17000 287200
rect 15800 284200 16000 284800
rect 16800 284200 17000 284800
rect 15800 281800 17000 284200
rect 15800 281200 16000 281800
rect 16800 281200 17000 281800
rect 15800 278800 17000 281200
rect 15800 278200 16000 278800
rect 16800 278200 17000 278800
rect 15800 275800 17000 278200
rect 15800 275200 16000 275800
rect 16800 275200 17000 275800
rect 15800 272800 17000 275200
rect 15800 272200 16000 272800
rect 16800 272200 17000 272800
rect 15800 269800 17000 272200
rect 15800 269200 16000 269800
rect 16800 269200 17000 269800
rect 15800 266800 17000 269200
rect 15800 266200 16000 266800
rect 16800 266200 17000 266800
rect 15800 263800 17000 266200
rect 15800 263200 16000 263800
rect 16800 263200 17000 263800
rect 15800 260800 17000 263200
rect 15800 260200 16000 260800
rect 16800 260200 17000 260800
rect 15800 257800 17000 260200
rect 15800 257200 16000 257800
rect 16800 257200 17000 257800
rect 15800 254800 17000 257200
rect 15800 254200 16000 254800
rect 16800 254200 17000 254800
rect 15800 251800 17000 254200
rect 15800 251200 16000 251800
rect 16800 251200 17000 251800
rect 15800 248800 17000 251200
rect 15800 248200 16000 248800
rect 16800 248200 17000 248800
rect 15800 245800 17000 248200
rect 15800 245200 16000 245800
rect 16800 245200 17000 245800
rect 15800 242800 17000 245200
rect 15800 242200 16000 242800
rect 16800 242200 17000 242800
rect 15800 239800 17000 242200
rect 15800 239200 16000 239800
rect 16800 239200 17000 239800
rect 15800 236800 17000 239200
rect 15800 236200 16000 236800
rect 16800 236200 17000 236800
rect 15800 233800 17000 236200
rect 15800 233200 16000 233800
rect 16800 233200 17000 233800
rect 15800 230800 17000 233200
rect 15800 230200 16000 230800
rect 16800 230200 17000 230800
rect 15800 227800 17000 230200
rect 15800 227200 16000 227800
rect 16800 227200 17000 227800
rect 15800 224800 17000 227200
rect 15800 224200 16000 224800
rect 16800 224200 17000 224800
rect 15800 221800 17000 224200
rect 15800 221200 16000 221800
rect 16800 221200 17000 221800
rect 15800 218800 17000 221200
rect 15800 218200 16000 218800
rect 16800 218200 17000 218800
rect 15800 215800 17000 218200
rect 15800 215200 16000 215800
rect 16800 215200 17000 215800
rect 15800 212800 17000 215200
rect 15800 212200 16000 212800
rect 16800 212200 17000 212800
rect 15800 209800 17000 212200
rect 15800 209200 16000 209800
rect 16800 209200 17000 209800
rect 15800 206800 17000 209200
rect 15800 206200 16000 206800
rect 16800 206200 17000 206800
rect 15800 203800 17000 206200
rect 15800 203200 16000 203800
rect 16800 203200 17000 203800
rect 15800 200800 17000 203200
rect 15800 200200 16000 200800
rect 16800 200200 17000 200800
rect 15800 197800 17000 200200
rect 15800 197200 16000 197800
rect 16800 197200 17000 197800
rect 15800 194800 17000 197200
rect 15800 194200 16000 194800
rect 16800 194200 17000 194800
rect 15800 191800 17000 194200
rect 15800 191200 16000 191800
rect 16800 191200 17000 191800
rect 15800 188800 17000 191200
rect 15800 188200 16000 188800
rect 16800 188200 17000 188800
rect 15800 185800 17000 188200
rect 15800 185200 16000 185800
rect 16800 185200 17000 185800
rect 15800 182800 17000 185200
rect 15800 182200 16000 182800
rect 16800 182200 17000 182800
rect 15800 179800 17000 182200
rect 15800 179200 16000 179800
rect 16800 179200 17000 179800
rect 400 177370 2740 177720
rect 400 163110 700 177370
rect 2330 163110 2740 177370
rect 400 162870 2740 163110
rect 15800 176800 17000 179200
rect 15800 176200 16000 176800
rect 16800 176200 17000 176800
rect 15800 173800 17000 176200
rect 15800 173200 16000 173800
rect 16800 173200 17000 173800
rect 15800 170800 17000 173200
rect 15800 170200 16000 170800
rect 16800 170200 17000 170800
rect 15800 167800 17000 170200
rect 15800 167200 16000 167800
rect 16800 167200 17000 167800
rect 15800 164800 17000 167200
rect 15800 164200 16000 164800
rect 16800 164200 17000 164800
rect 15800 161800 17000 164200
rect 15800 161200 16000 161800
rect 16800 161200 17000 161800
rect 15800 158800 17000 161200
rect 15800 158200 16000 158800
rect 16800 158200 17000 158800
rect 15800 155800 17000 158200
rect 15800 155200 16000 155800
rect 16800 155200 17000 155800
rect 15800 152800 17000 155200
rect 15800 152200 16000 152800
rect 16800 152200 17000 152800
rect 15800 149800 17000 152200
rect 15800 149200 16000 149800
rect 16800 149200 17000 149800
rect 15800 146800 17000 149200
rect 15800 146200 16000 146800
rect 16800 146200 17000 146800
rect 15800 143800 17000 146200
rect 15800 143200 16000 143800
rect 16800 143200 17000 143800
rect 15800 140800 17000 143200
rect 15800 140200 16000 140800
rect 16800 140200 17000 140800
rect 15800 137800 17000 140200
rect 15800 137200 16000 137800
rect 16800 137200 17000 137800
rect 15800 134800 17000 137200
rect 15800 134200 16000 134800
rect 16800 134200 17000 134800
rect 15800 131800 17000 134200
rect 15800 131200 16000 131800
rect 16800 131200 17000 131800
rect 15800 128800 17000 131200
rect 15800 128200 16000 128800
rect 16800 128200 17000 128800
rect 15800 125800 17000 128200
rect 15800 125200 16000 125800
rect 16800 125200 17000 125800
rect 15800 122800 17000 125200
rect 15800 122200 16000 122800
rect 16800 122200 17000 122800
rect 15800 119800 17000 122200
rect 15800 119200 16000 119800
rect 16800 119200 17000 119800
rect 15800 116800 17000 119200
rect 15800 116200 16000 116800
rect 16800 116200 17000 116800
rect 15800 113800 17000 116200
rect 15800 113200 16000 113800
rect 16800 113200 17000 113800
rect 15800 110800 17000 113200
rect 15800 110200 16000 110800
rect 16800 110200 17000 110800
rect 15800 107800 17000 110200
rect 15800 107200 16000 107800
rect 16800 107200 17000 107800
rect 15800 104800 17000 107200
rect 15800 104200 16000 104800
rect 16800 104200 17000 104800
rect 15800 101800 17000 104200
rect 15800 101200 16000 101800
rect 16800 101200 17000 101800
rect 15800 98800 17000 101200
rect 15800 98200 16000 98800
rect 16800 98200 17000 98800
rect 15800 95800 17000 98200
rect 15800 95200 16000 95800
rect 16800 95200 17000 95800
rect 15800 92800 17000 95200
rect 15800 92200 16000 92800
rect 16800 92200 17000 92800
rect 15800 89800 17000 92200
rect 15800 89200 16000 89800
rect 16800 89200 17000 89800
rect 15800 86800 17000 89200
rect 15800 86200 16000 86800
rect 16800 86200 17000 86800
rect 15800 83800 17000 86200
rect 15800 83200 16000 83800
rect 16800 83200 17000 83800
rect 15800 80800 17000 83200
rect 15800 80200 16000 80800
rect 16800 80200 17000 80800
rect 15800 77800 17000 80200
rect 15800 77200 16000 77800
rect 16800 77200 17000 77800
rect 15800 74800 17000 77200
rect 15800 74200 16000 74800
rect 16800 74200 17000 74800
rect 15800 71800 17000 74200
rect 15800 71200 16000 71800
rect 16800 71200 17000 71800
rect 15800 68800 17000 71200
rect 15800 68200 16000 68800
rect 16800 68200 17000 68800
rect 15800 65800 17000 68200
rect 15800 65200 16000 65800
rect 16800 65200 17000 65800
rect 15800 62800 17000 65200
rect 15800 62200 16000 62800
rect 16800 62200 17000 62800
rect 15800 59800 17000 62200
rect 15800 59200 16000 59800
rect 16800 59200 17000 59800
rect 15800 56800 17000 59200
rect 15800 56200 16000 56800
rect 16800 56200 17000 56800
rect 15800 53800 17000 56200
rect 15800 53200 16000 53800
rect 16800 53200 17000 53800
rect 15800 50800 17000 53200
rect 15800 50200 16000 50800
rect 16800 50200 17000 50800
rect 15800 47800 17000 50200
rect 15800 47200 16000 47800
rect 16800 47200 17000 47800
rect 15800 44800 17000 47200
rect 15800 44200 16000 44800
rect 16800 44200 17000 44800
rect 15800 41800 17000 44200
rect 15800 41200 16000 41800
rect 16800 41200 17000 41800
rect 15800 38800 17000 41200
rect 15800 38200 16000 38800
rect 16800 38200 17000 38800
rect 15800 35800 17000 38200
rect 15800 35200 16000 35800
rect 16800 35200 17000 35800
rect 15800 32800 17000 35200
rect 15800 32200 16000 32800
rect 16800 32200 17000 32800
rect 15800 29800 17000 32200
rect 15800 29200 16000 29800
rect 16800 29200 17000 29800
rect 15800 26800 17000 29200
rect 15800 26200 16000 26800
rect 16800 26200 17000 26800
rect 15800 23800 17000 26200
rect 15800 23200 16000 23800
rect 16800 23200 17000 23800
rect 15800 20800 17000 23200
rect 15800 20200 16000 20800
rect 16800 20200 17000 20800
rect 15800 17800 17000 20200
rect 15800 17200 16000 17800
rect 16800 17200 17000 17800
rect 15800 14800 17000 17200
rect 15800 14200 16000 14800
rect 16800 14200 17000 14800
rect 15800 11800 17000 14200
rect 15800 11200 16000 11800
rect 16800 11200 17000 11800
rect 15800 8800 17000 11200
rect 15800 8200 16000 8800
rect 16800 8200 17000 8800
rect 15800 5800 17000 8200
rect 15800 5200 16000 5800
rect 16800 5200 17000 5800
rect 15800 4400 17000 5200
rect 475200 330000 475800 331400
rect 477200 330000 477800 331400
rect 475200 329400 477800 330000
rect 475200 328000 475800 329400
rect 477200 328000 477800 329400
rect 475200 327400 477800 328000
rect 475200 326000 475800 327400
rect 477200 326000 477800 327400
rect 475200 325400 477800 326000
rect 475200 324000 475800 325400
rect 477200 324000 477800 325400
rect 475200 323400 477800 324000
rect 475200 322000 475800 323400
rect 477200 322000 477800 323400
rect 475200 321400 477800 322000
rect 475200 320000 475800 321400
rect 477200 320000 477800 321400
rect 475200 319400 477800 320000
rect 475200 318000 475800 319400
rect 477200 318000 477800 319400
rect 475200 317400 477800 318000
rect 475200 316000 475800 317400
rect 477200 316000 477800 317400
rect 475200 315400 477800 316000
rect 475200 314000 475800 315400
rect 477200 314000 477800 315400
rect 475200 313400 477800 314000
rect 475200 312000 475800 313400
rect 477200 312000 477800 313400
rect 475200 311400 477800 312000
rect 475200 310000 475800 311400
rect 477200 310000 477800 311400
rect 475200 309400 477800 310000
rect 475200 308000 475800 309400
rect 477200 308000 477800 309400
rect 475200 307400 477800 308000
rect 475200 306000 475800 307400
rect 477200 306000 477800 307400
rect 475200 305400 477800 306000
rect 475200 304000 475800 305400
rect 477200 304000 477800 305400
rect 475200 303400 477800 304000
rect 475200 302000 475800 303400
rect 477200 302000 477800 303400
rect 475200 301400 477800 302000
rect 475200 300000 475800 301400
rect 477200 300000 477800 301400
rect 475200 299400 477800 300000
rect 475200 298000 475800 299400
rect 477200 298000 477800 299400
rect 475200 297400 477800 298000
rect 475200 296000 475800 297400
rect 477200 296000 477800 297400
rect 475200 295400 477800 296000
rect 475200 294000 475800 295400
rect 477200 294000 477800 295400
rect 475200 293400 477800 294000
rect 475200 292000 475800 293400
rect 477200 292000 477800 293400
rect 475200 291400 477800 292000
rect 475200 290000 475800 291400
rect 477200 290000 477800 291400
rect 475200 289400 477800 290000
rect 475200 288000 475800 289400
rect 477200 288000 477800 289400
rect 475200 287400 477800 288000
rect 475200 286000 475800 287400
rect 477200 286000 477800 287400
rect 475200 285400 477800 286000
rect 475200 284000 475800 285400
rect 477200 284000 477800 285400
rect 475200 283400 477800 284000
rect 475200 282000 475800 283400
rect 477200 282000 477800 283400
rect 475200 281400 477800 282000
rect 475200 280000 475800 281400
rect 477200 280000 477800 281400
rect 475200 279400 477800 280000
rect 475200 278000 475800 279400
rect 477200 278000 477800 279400
rect 475200 277400 477800 278000
rect 475200 276000 475800 277400
rect 477200 276000 477800 277400
rect 475200 275400 477800 276000
rect 475200 274000 475800 275400
rect 477200 274000 477800 275400
rect 475200 273400 477800 274000
rect 475200 272000 475800 273400
rect 477200 272000 477800 273400
rect 475200 271400 477800 272000
rect 475200 270000 475800 271400
rect 477200 270000 477800 271400
rect 475200 269400 477800 270000
rect 475200 268000 475800 269400
rect 477200 268000 477800 269400
rect 475200 267400 477800 268000
rect 475200 266000 475800 267400
rect 477200 266000 477800 267400
rect 475200 265400 477800 266000
rect 475200 264000 475800 265400
rect 477200 264000 477800 265400
rect 475200 263400 477800 264000
rect 475200 262000 475800 263400
rect 477200 262000 477800 263400
rect 475200 261400 477800 262000
rect 475200 260000 475800 261400
rect 477200 260000 477800 261400
rect 475200 259400 477800 260000
rect 475200 258000 475800 259400
rect 477200 258000 477800 259400
rect 568800 453000 582400 468600
rect 568800 366400 573400 453000
rect 576400 396400 582600 397600
rect 576400 395800 576800 396400
rect 582200 395800 582600 396400
rect 576400 394400 582600 395800
rect 576400 393800 576800 394400
rect 582200 393800 582600 394400
rect 576400 392400 582600 393800
rect 576400 391800 576800 392400
rect 582200 391800 582600 392400
rect 576400 390400 582600 391800
rect 576400 389800 576800 390400
rect 582200 389800 582600 390400
rect 576400 388400 582600 389800
rect 576400 387800 576800 388400
rect 582200 387800 582600 388400
rect 576400 386400 582600 387800
rect 576400 385800 576800 386400
rect 582200 385800 582600 386400
rect 576400 384400 582600 385800
rect 576400 383800 576800 384400
rect 582200 383800 582600 384400
rect 576400 382400 582600 383800
rect 576400 381800 576800 382400
rect 582200 381800 582600 382400
rect 576400 380400 582600 381800
rect 576400 379800 576800 380400
rect 582200 379800 582600 380400
rect 576400 378400 582600 379800
rect 576400 377800 576800 378400
rect 582200 377800 582600 378400
rect 576400 376400 582600 377800
rect 576400 375800 576800 376400
rect 582200 375800 582600 376400
rect 576400 374400 582600 375800
rect 576400 373800 576800 374400
rect 582200 373800 582600 374400
rect 576400 372400 582600 373800
rect 576400 371800 576800 372400
rect 582200 371800 582600 372400
rect 576400 370400 582600 371800
rect 576400 369800 576800 370400
rect 582200 369800 582600 370400
rect 576400 369400 582600 369800
rect 568800 365400 579200 366400
rect 568800 361800 573400 365400
rect 573800 364800 574800 365200
rect 573800 363400 574000 364800
rect 574600 363400 574800 364800
rect 573800 363000 574800 363400
rect 575600 365000 576400 365400
rect 575600 363400 575800 365000
rect 576000 363400 576400 365000
rect 575600 363200 576400 363400
rect 576600 364800 577600 365200
rect 576600 363400 576800 364800
rect 577400 363400 577600 364800
rect 576600 363000 577600 363400
rect 578400 365000 579200 365400
rect 578400 363400 578600 365000
rect 578800 363400 579200 365000
rect 578400 363200 579200 363400
rect 579600 363000 582400 369400
rect 573800 362400 582400 363000
rect 568800 361400 574800 361800
rect 577360 361700 582400 362400
rect 568800 361200 572600 361400
rect 573400 361200 573800 361400
rect 574600 361200 574800 361400
rect 568800 361000 574800 361200
rect 568800 360800 572600 361000
rect 573400 360800 573800 361000
rect 574600 360800 574800 361000
rect 568800 360600 574800 360800
rect 568800 360400 572600 360600
rect 573400 360400 573800 360600
rect 574600 360400 574800 360600
rect 568800 360200 574800 360400
rect 568800 360000 572600 360200
rect 573400 360000 573800 360200
rect 574600 360000 574800 360200
rect 568800 359800 574800 360000
rect 568800 359600 572600 359800
rect 573400 359600 573800 359800
rect 574600 359600 574800 359800
rect 568800 359400 574800 359600
rect 568800 359200 572600 359400
rect 573400 359200 573800 359400
rect 574600 359200 574800 359400
rect 568800 359000 574800 359200
rect 568800 358800 572600 359000
rect 573400 358800 573800 359000
rect 574600 358800 574800 359000
rect 568800 358600 574800 358800
rect 568800 358400 572600 358600
rect 573400 358400 573800 358600
rect 574600 358400 574800 358600
rect 568800 358200 574800 358400
rect 568800 358000 572600 358200
rect 573400 358000 573800 358200
rect 574600 358000 574800 358200
rect 568800 357800 574800 358000
rect 568800 357600 572600 357800
rect 573400 357600 573800 357800
rect 574600 357600 574800 357800
rect 568800 357400 574800 357600
rect 568800 357200 572600 357400
rect 573400 357200 573800 357400
rect 574600 357200 574800 357400
rect 568800 357000 574800 357200
rect 568800 356800 572600 357000
rect 573400 356800 573800 357000
rect 574600 356800 574800 357000
rect 568800 356600 574800 356800
rect 577420 361200 582400 361700
rect 577420 356720 578780 361200
rect 568800 356400 572600 356600
rect 573400 356400 573800 356600
rect 574600 356400 574800 356600
rect 568800 356200 574800 356400
rect 568800 356000 572600 356200
rect 573400 356000 573800 356200
rect 574600 356000 574800 356200
rect 568800 355800 574800 356000
rect 568800 355600 572600 355800
rect 573400 355600 573800 355800
rect 574600 355600 574800 355800
rect 568800 355400 574800 355600
rect 568800 355200 572600 355400
rect 573400 355200 573800 355400
rect 574600 355200 574800 355400
rect 568800 355000 574800 355200
rect 568800 354800 572600 355000
rect 573400 354800 573800 355000
rect 574600 354800 574800 355000
rect 568800 354600 574800 354800
rect 568800 354400 572600 354600
rect 573400 354400 573800 354600
rect 574600 354400 574800 354600
rect 577410 356710 581180 356720
rect 577410 354570 582860 356710
rect 568800 354200 574800 354400
rect 568800 354000 572600 354200
rect 573400 354000 573800 354200
rect 574600 354000 574800 354200
rect 568800 353800 574800 354000
rect 568800 271600 572000 353800
rect 568800 270600 569200 271600
rect 571600 270600 572000 271600
rect 568800 269600 572000 270600
rect 568800 268600 569200 269600
rect 571600 268600 572000 269600
rect 568800 267600 572000 268600
rect 568800 266600 569200 267600
rect 571600 266600 572000 267600
rect 568800 265600 572000 266600
rect 580840 266510 582860 354570
rect 568800 264600 569200 265600
rect 571600 264600 572000 265600
rect 568800 263600 572000 264600
rect 568800 262600 569200 263600
rect 571600 262600 572000 263600
rect 568800 261600 572000 262600
rect 568800 260600 569200 261600
rect 571600 260600 572000 261600
rect 568800 259600 572000 260600
rect 568800 258600 569200 259600
rect 571600 258600 572000 259600
rect 568800 258200 572000 258600
rect 580430 265330 583850 266510
rect 580430 264550 580810 265330
rect 583470 264550 583850 265330
rect 580430 263500 583850 264550
rect 580430 262720 580840 263500
rect 583500 262720 583850 263500
rect 580430 261910 583850 262720
rect 580430 261130 580810 261910
rect 583470 261130 583850 261910
rect 580430 260290 583850 261130
rect 580430 259510 580780 260290
rect 583440 259510 583850 260290
rect 580430 259100 583850 259510
rect 580430 258320 580810 259100
rect 583470 258320 583850 259100
rect 475200 257400 477800 258000
rect 580430 257890 583850 258320
rect 475200 256000 475800 257400
rect 477200 256000 477800 257400
rect 475200 255400 477800 256000
rect 475200 254000 475800 255400
rect 477200 254000 477800 255400
rect 475200 253400 477800 254000
rect 475200 252000 475800 253400
rect 477200 252000 477800 253400
rect 475200 251400 477800 252000
rect 475200 250000 475800 251400
rect 477200 250000 477800 251400
rect 475200 249400 477800 250000
rect 475200 248000 475800 249400
rect 477200 248000 477800 249400
rect 475200 247400 477800 248000
rect 475200 246000 475800 247400
rect 477200 246000 477800 247400
rect 475200 245400 477800 246000
rect 475200 244000 475800 245400
rect 477200 244000 477800 245400
rect 475200 243400 477800 244000
rect 475200 242000 475800 243400
rect 477200 242000 477800 243400
rect 475200 241400 477800 242000
rect 475200 240000 475800 241400
rect 477200 240000 477800 241400
rect 568600 241530 577600 242800
rect 568600 240370 568700 241530
rect 569770 241520 577600 241530
rect 577420 240400 577600 241520
rect 576370 240370 577600 240400
rect 568600 240310 577600 240370
rect 475200 239400 477800 240000
rect 475200 238000 475800 239400
rect 477200 238000 477800 239400
rect 475200 237400 477800 238000
rect 475200 236000 475800 237400
rect 477200 236000 477800 237400
rect 475200 235400 477800 236000
rect 475200 234000 475800 235400
rect 477200 234000 477800 235400
rect 475200 233400 477800 234000
rect 475200 232000 475800 233400
rect 477200 232000 477800 233400
rect 475200 231400 477800 232000
rect 475200 230000 475800 231400
rect 477200 230000 477800 231400
rect 475200 229400 477800 230000
rect 475200 228000 475800 229400
rect 477200 228000 477800 229400
rect 475200 227400 477800 228000
rect 475200 226000 475800 227400
rect 477200 226000 477800 227400
rect 475200 225400 477800 226000
rect 475200 224000 475800 225400
rect 477200 224000 477800 225400
rect 475200 223400 477800 224000
rect 475200 222000 475800 223400
rect 477200 222000 477800 223400
rect 475200 221400 477800 222000
rect 475200 220000 475800 221400
rect 477200 220000 477800 221400
rect 475200 219400 477800 220000
rect 475200 218000 475800 219400
rect 477200 218000 477800 219400
rect 475200 217400 477800 218000
rect 475200 216000 475800 217400
rect 477200 216000 477800 217400
rect 567650 240000 577600 240310
rect 567650 239920 572500 240000
rect 567650 217220 568050 239920
rect 572020 217610 572260 217640
rect 572020 217220 572040 217610
rect 567650 216820 572040 217220
rect 572020 216420 572040 216820
rect 572230 216420 572260 217610
rect 572020 216390 572260 216420
rect 475200 215400 477800 216000
rect 475200 214000 475800 215400
rect 477200 214000 477800 215400
rect 475200 213400 477800 214000
rect 475200 212000 475800 213400
rect 477200 212000 477800 213400
rect 475200 211400 477800 212000
rect 475200 210000 475800 211400
rect 477200 210000 477800 211400
rect 475200 209400 477800 210000
rect 475200 208000 475800 209400
rect 477200 208000 477800 209400
rect 475200 207400 477800 208000
rect 475200 206000 475800 207400
rect 477200 206000 477800 207400
rect 475200 205400 477800 206000
rect 475200 204000 475800 205400
rect 477200 204000 477800 205400
rect 475200 203400 477800 204000
rect 475200 202000 475800 203400
rect 477200 202000 477800 203400
rect 475200 201400 477800 202000
rect 475200 200000 475800 201400
rect 477200 200000 477800 201400
rect 475200 199400 477800 200000
rect 475200 198000 475800 199400
rect 477200 198000 477800 199400
rect 475200 197400 477800 198000
rect 475200 196000 475800 197400
rect 477200 196000 477800 197400
rect 475200 195400 477800 196000
rect 475200 194000 475800 195400
rect 477200 194000 477800 195400
rect 475200 193400 477800 194000
rect 475200 192000 475800 193400
rect 477200 192000 477800 193400
rect 475200 191400 477800 192000
rect 475200 190000 475800 191400
rect 477200 190000 477800 191400
rect 475200 189400 477800 190000
rect 579200 201000 581200 201200
rect 579200 198160 579460 201000
rect 580960 198160 581200 201000
rect 579200 189900 579500 198160
rect 580900 189900 581200 198160
rect 579200 189500 581200 189900
rect 475200 188000 475800 189400
rect 477200 188000 477800 189400
rect 475200 187400 477800 188000
rect 475200 186000 475800 187400
rect 477200 186000 477800 187400
rect 475200 185400 477800 186000
rect 475200 184000 475800 185400
rect 477200 184000 477800 185400
rect 475200 183400 477800 184000
rect 475200 182000 475800 183400
rect 477200 182000 477800 183400
rect 475200 181400 477800 182000
rect 475200 180000 475800 181400
rect 477200 180000 477800 181400
rect 475200 179400 477800 180000
rect 475200 178000 475800 179400
rect 477200 178000 477800 179400
rect 475200 177400 477800 178000
rect 475200 176000 475800 177400
rect 477200 176000 477800 177400
rect 475200 175400 477800 176000
rect 475200 174000 475800 175400
rect 477200 174000 477800 175400
rect 475200 173400 477800 174000
rect 475200 172000 475800 173400
rect 477200 172000 477800 173400
rect 475200 171400 477800 172000
rect 475200 170000 475800 171400
rect 477200 170000 477800 171400
rect 475200 169400 477800 170000
rect 475200 168000 475800 169400
rect 477200 168000 477800 169400
rect 475200 167400 477800 168000
rect 475200 166000 475800 167400
rect 477200 166000 477800 167400
rect 576200 175500 579600 175800
rect 576200 167200 576400 175500
rect 579400 167200 579600 175500
rect 576200 166600 579600 167200
rect 475200 165400 477800 166000
rect 475200 164000 475800 165400
rect 477200 164000 477800 165400
rect 475200 163400 477800 164000
rect 475200 162000 475800 163400
rect 477200 162000 477800 163400
rect 475200 161400 477800 162000
rect 475200 160000 475800 161400
rect 477200 160000 477800 161400
rect 475200 159400 477800 160000
rect 475200 158000 475800 159400
rect 477200 158000 477800 159400
rect 475200 157400 477800 158000
rect 475200 156000 475800 157400
rect 477200 156000 477800 157400
rect 475200 155400 477800 156000
rect 475200 154000 475800 155400
rect 477200 154000 477800 155400
rect 475200 153400 477800 154000
rect 475200 152000 475800 153400
rect 477200 152000 477800 153400
rect 475200 151400 477800 152000
rect 475200 150000 475800 151400
rect 477200 150000 477800 151400
rect 475200 149400 477800 150000
rect 475200 148000 475800 149400
rect 477200 148000 477800 149400
rect 475200 147400 477800 148000
rect 475200 146000 475800 147400
rect 477200 146000 477800 147400
rect 475200 145400 477800 146000
rect 475200 144000 475800 145400
rect 477200 144000 477800 145400
rect 475200 143400 477800 144000
rect 475200 142000 475800 143400
rect 477200 142000 477800 143400
rect 572900 152000 576700 152600
rect 572900 151830 573200 152000
rect 572900 148990 573150 151830
rect 572900 143700 573200 148990
rect 576200 143700 576700 152000
rect 572900 143300 576700 143700
rect 475200 141400 477800 142000
rect 475200 140000 475800 141400
rect 477200 140000 477800 141400
rect 475200 139400 477800 140000
rect 475200 138000 475800 139400
rect 477200 138000 477800 139400
rect 475200 137400 477800 138000
rect 475200 136000 475800 137400
rect 477200 136000 477800 137400
rect 475200 135400 477800 136000
rect 475200 134000 475800 135400
rect 477200 134000 477800 135400
rect 475200 133400 477800 134000
rect 475200 132000 475800 133400
rect 477200 132000 477800 133400
rect 475200 131400 477800 132000
rect 475200 130000 475800 131400
rect 477200 130000 477800 131400
rect 475200 129400 477800 130000
rect 475200 128000 475800 129400
rect 477200 128000 477800 129400
rect 475200 127400 477800 128000
rect 475200 126000 475800 127400
rect 477200 126000 477800 127400
rect 475200 125400 477800 126000
rect 475200 124000 475800 125400
rect 477200 124000 477800 125400
rect 475200 123400 477800 124000
rect 475200 122000 475800 123400
rect 477200 122000 477800 123400
rect 570290 130870 578040 131480
rect 570290 130770 570900 130870
rect 570290 123400 570850 130770
rect 577350 123430 578040 130870
rect 577320 123400 578040 123430
rect 570290 123020 578040 123400
rect 475200 121400 477800 122000
rect 475200 120000 475800 121400
rect 477200 120000 477800 121400
rect 475200 119400 477800 120000
rect 475200 118000 475800 119400
rect 477200 118000 477800 119400
rect 475200 117400 477800 118000
rect 475200 116000 475800 117400
rect 477200 116000 477800 117400
rect 475200 115400 477800 116000
rect 475200 114000 475800 115400
rect 477200 114000 477800 115400
rect 475200 113400 477800 114000
rect 475200 112000 475800 113400
rect 477200 112000 477800 113400
rect 475200 111400 477800 112000
rect 475200 110000 475800 111400
rect 477200 110000 477800 111400
rect 475200 109400 477800 110000
rect 475200 108000 475800 109400
rect 477200 108000 477800 109400
rect 475200 107400 477800 108000
rect 475200 106000 475800 107400
rect 477200 106000 477800 107400
rect 475200 105400 477800 106000
rect 475200 104000 475800 105400
rect 477200 104000 477800 105400
rect 475200 103400 477800 104000
rect 475200 102000 475800 103400
rect 477200 102000 477800 103400
rect 475200 101400 477800 102000
rect 475200 100000 475800 101400
rect 477200 100000 477800 101400
rect 475200 99400 477800 100000
rect 475200 98000 475800 99400
rect 477200 98000 477800 99400
rect 475200 97400 477800 98000
rect 475200 96000 475800 97400
rect 477200 96000 477800 97400
rect 475200 95400 477800 96000
rect 475200 94000 475800 95400
rect 477200 94000 477800 95400
rect 475200 93400 477800 94000
rect 475200 92000 475800 93400
rect 477200 92000 477800 93400
rect 475200 91400 477800 92000
rect 475200 90000 475800 91400
rect 477200 90000 477800 91400
rect 475200 89400 477800 90000
rect 475200 88000 475800 89400
rect 477200 88000 477800 89400
rect 475200 87400 477800 88000
rect 475200 86000 475800 87400
rect 477200 86000 477800 87400
rect 475200 85400 477800 86000
rect 475200 84000 475800 85400
rect 477200 84000 477800 85400
rect 475200 83400 477800 84000
rect 475200 82000 475800 83400
rect 477200 82000 477800 83400
rect 475200 81400 477800 82000
rect 475200 80000 475800 81400
rect 477200 80000 477800 81400
rect 475200 79400 477800 80000
rect 475200 78000 475800 79400
rect 477200 78000 477800 79400
rect 475200 77400 477800 78000
rect 475200 76000 475800 77400
rect 477200 76000 477800 77400
rect 475200 75400 477800 76000
rect 475200 74000 475800 75400
rect 477200 74000 477800 75400
rect 475200 73400 477800 74000
rect 475200 72000 475800 73400
rect 477200 72000 477800 73400
rect 475200 71400 477800 72000
rect 475200 70000 475800 71400
rect 477200 70000 477800 71400
rect 475200 69400 477800 70000
rect 475200 68000 475800 69400
rect 477200 68000 477800 69400
rect 475200 67400 477800 68000
rect 475200 66000 475800 67400
rect 477200 66000 477800 67400
rect 475200 65400 477800 66000
rect 475200 64000 475800 65400
rect 477200 64000 477800 65400
rect 475200 63400 477800 64000
rect 475200 62000 475800 63400
rect 477200 62000 477800 63400
rect 475200 61400 477800 62000
rect 475200 60000 475800 61400
rect 477200 60000 477800 61400
rect 475200 59400 477800 60000
rect 475200 58000 475800 59400
rect 477200 58000 477800 59400
rect 475200 57400 477800 58000
rect 475200 56000 475800 57400
rect 477200 56000 477800 57400
rect 475200 55400 477800 56000
rect 475200 54000 475800 55400
rect 477200 54000 477800 55400
rect 475200 53400 477800 54000
rect 475200 52000 475800 53400
rect 477200 52000 477800 53400
rect 475200 51400 477800 52000
rect 475200 50000 475800 51400
rect 477200 50000 477800 51400
rect 475200 49400 477800 50000
rect 475200 48000 475800 49400
rect 477200 48000 477800 49400
rect 475200 47400 477800 48000
rect 475200 46000 475800 47400
rect 477200 46000 477800 47400
rect 475200 45400 477800 46000
rect 475200 44000 475800 45400
rect 477200 44000 477800 45400
rect 475200 43400 477800 44000
rect 475200 42000 475800 43400
rect 477200 42000 477800 43400
rect 475200 41400 477800 42000
rect 475200 40000 475800 41400
rect 477200 40000 477800 41400
rect 475200 39400 477800 40000
rect 475200 38000 475800 39400
rect 477200 38000 477800 39400
rect 475200 37400 477800 38000
rect 475200 36000 475800 37400
rect 477200 36000 477800 37400
rect 475200 35400 477800 36000
rect 475200 34000 475800 35400
rect 477200 34000 477800 35400
rect 475200 33400 477800 34000
rect 475200 32000 475800 33400
rect 477200 32000 477800 33400
rect 475200 31400 477800 32000
rect 475200 30000 475800 31400
rect 477200 30000 477800 31400
rect 475200 29400 477800 30000
rect 475200 28000 475800 29400
rect 477200 28000 477800 29400
rect 475200 27400 477800 28000
rect 475200 26000 475800 27400
rect 477200 26000 477800 27400
rect 475200 25400 477800 26000
rect 475200 24000 475800 25400
rect 477200 24000 477800 25400
rect 475200 23400 477800 24000
rect 475200 22000 475800 23400
rect 477200 22000 477800 23400
rect 475200 21400 477800 22000
rect 475200 20000 475800 21400
rect 477200 20000 477800 21400
rect 475200 19400 477800 20000
rect 475200 18000 475800 19400
rect 477200 18000 477800 19400
rect 475200 17400 477800 18000
rect 475200 16000 475800 17400
rect 477200 16000 477800 17400
rect 475200 15400 477800 16000
rect 475200 14000 475800 15400
rect 477200 14000 477800 15400
rect 475200 13400 477800 14000
rect 475200 12000 475800 13400
rect 477200 12000 477800 13400
rect 475200 11400 477800 12000
rect 475200 10000 475800 11400
rect 477200 10000 477800 11400
rect 475200 9400 477800 10000
rect 475200 8000 475800 9400
rect 477200 8000 477800 9400
rect 475200 7400 477800 8000
rect 475200 6000 475800 7400
rect 477200 6000 477800 7400
rect 475200 5400 477800 6000
rect 475200 4400 475800 5400
rect 15800 4000 475800 4400
rect 477200 4400 477800 5400
rect 477200 4000 568600 4400
rect 15800 2200 568600 4000
rect 475200 2000 477800 2200
<< via4 >>
rect 228670 701850 232530 702520
rect 330480 701740 334340 702410
rect 222600 698000 226600 698800
rect 222600 696800 226600 697600
rect 222600 695600 226600 696400
rect 324200 698000 328200 698800
rect 324200 696800 328200 697600
rect 324200 695600 328200 696400
rect 510880 696600 525130 703440
rect 7200 690200 9000 691600
rect 11000 690200 12800 691600
rect 15800 690200 16800 691400
rect 18800 690200 19800 691400
rect 21800 690200 22800 691400
rect 24800 690200 25800 691400
rect 27800 690200 28800 691400
rect 30800 690200 31800 691400
rect 33800 690200 34800 691400
rect 36800 690200 37800 691400
rect 39800 690200 40800 691400
rect 42800 690200 43800 691400
rect 45800 690200 46800 691400
rect 48800 690200 49800 691400
rect 51800 690200 52800 691400
rect 54800 690200 55800 691400
rect 57800 690200 58800 691400
rect 60800 690200 61800 691400
rect 63800 690200 64800 691400
rect 66800 690200 67800 691400
rect 69800 690200 70800 691400
rect 72800 690200 73800 691400
rect 75800 690200 76800 691400
rect 78800 690200 79800 691400
rect 81800 690200 82800 691400
rect 84800 690200 85800 691400
rect 87800 690200 88800 691400
rect 90800 690200 91800 691400
rect 93800 690200 94800 691400
rect 96800 690200 97800 691400
rect 99800 690200 100800 691400
rect 102800 690200 103800 691400
rect 105800 690200 106800 691400
rect 108800 690200 109800 691400
rect 111800 690200 112800 691400
rect 114800 690200 115800 691400
rect 117800 690200 118800 691400
rect 120800 690200 121800 691400
rect 123800 690200 124800 691400
rect 126800 690200 127800 691400
rect 129800 690200 130800 691400
rect 132800 690200 133800 691400
rect 135800 690200 136800 691400
rect 138800 690200 139800 691400
rect 141800 690200 142800 691400
rect 144800 690200 145800 691400
rect 147800 690200 148800 691400
rect 150800 690200 151800 691400
rect 153800 690200 154800 691400
rect 156800 690200 157800 691400
rect 159800 690200 160800 691400
rect 162800 690200 163800 691400
rect 165800 690200 166800 691400
rect 168800 690200 169800 691400
rect 171800 690200 172800 691400
rect 174800 690200 175800 691400
rect 177800 690200 178800 691400
rect 180800 690200 181800 691400
rect 183800 690200 184800 691400
rect 186800 690200 187800 691400
rect 189800 690200 190800 691400
rect 192800 690200 193800 691400
rect 195800 690200 196800 691400
rect 198800 690200 199800 691400
rect 201800 690200 202800 691400
rect 204800 690200 205800 691400
rect 207800 690200 208800 691400
rect 210800 690200 211800 691400
rect 213800 690200 214800 691400
rect 216800 690200 217800 691400
rect 219800 690200 220800 691400
rect 222800 690200 223800 691400
rect 225800 690200 226800 691400
rect 228800 690200 229800 691400
rect 231800 690200 232800 691400
rect 234800 690200 235800 691400
rect 237800 690200 238800 691400
rect 240800 690200 241800 691400
rect 243800 690200 244800 691400
rect 246800 690200 247800 691400
rect 249800 690200 250800 691400
rect 252800 690200 253800 691400
rect 255800 690200 256800 691400
rect 258800 690200 259800 691400
rect 261800 690200 262800 691400
rect 264800 690200 265800 691400
rect 267800 690200 268800 691400
rect 270800 690200 271800 691400
rect 273800 690200 274800 691400
rect 276800 690200 277800 691400
rect 279800 690200 280800 691400
rect 282800 690200 283800 691400
rect 285800 690200 286800 691400
rect 288800 690200 289800 691400
rect 291800 690200 292800 691400
rect 294800 690200 295800 691400
rect 297800 690200 298800 691400
rect 300800 690200 301800 691400
rect 303800 690200 304800 691400
rect 306800 690200 307800 691400
rect 309800 690200 310800 691400
rect 312800 690200 313800 691400
rect 315800 690200 316800 691400
rect 318800 690200 319800 691400
rect 321800 690200 322800 691400
rect 324800 690200 325800 691400
rect 327800 690200 328800 691400
rect 330800 690200 331800 691400
rect 333800 690200 334800 691400
rect 336800 690200 337800 691400
rect 339800 690200 340800 691400
rect 342800 690200 343800 691400
rect 345800 690200 346800 691400
rect 348800 690200 349800 691400
rect 351800 690200 352800 691400
rect 354800 690200 355800 691400
rect 357800 690200 358800 691400
rect 360800 690200 361800 691400
rect 363800 690200 364800 691400
rect 366800 690200 367800 691400
rect 369800 690200 370800 691400
rect 372800 690200 373800 691400
rect 375800 690200 376800 691400
rect 378800 690200 379800 691400
rect 381800 690200 382800 691400
rect 384800 690200 385800 691400
rect 387800 690200 388800 691400
rect 390800 690200 391800 691400
rect 393800 690200 394800 691400
rect 396800 690200 397800 691400
rect 399800 690200 400800 691400
rect 402800 690200 403800 691400
rect 405800 690200 406800 691400
rect 408800 690200 409800 691400
rect 411800 690200 412800 691400
rect 414800 690200 415800 691400
rect 417800 690200 418800 691400
rect 420800 690200 421800 691400
rect 423800 690200 424800 691400
rect 426800 690200 427800 691400
rect 429800 690200 430800 691400
rect 432800 690200 433800 691400
rect 435800 690200 436800 691400
rect 438800 690200 439800 691400
rect 441800 690200 442800 691400
rect 444800 690200 445800 691400
rect 447800 690200 448800 691400
rect 450800 690200 451800 691400
rect 453800 690200 454800 691400
rect 456800 690200 457800 691400
rect 459800 690200 460800 691400
rect 462800 690200 463800 691400
rect 465800 690200 466800 691400
rect 468800 690200 469800 691400
rect 471800 690200 472800 691400
rect 474800 690200 475800 691400
rect 477800 690200 478800 691400
rect 480800 690200 481800 691400
rect 483800 690200 484800 691400
rect 486800 690200 487800 691400
rect 489800 690200 490800 691400
rect 492800 690200 493800 691400
rect 495800 690200 496800 691400
rect 498800 690200 499800 691400
rect 501800 690200 502800 691400
rect 504800 690200 505800 691400
rect 507800 690200 508800 691400
rect 510800 690200 511800 691400
rect 513800 690200 514800 691400
rect 516800 690200 517800 691400
rect 519800 690200 520800 691400
rect 522800 690200 523800 691400
rect 525800 690200 526800 691400
rect 528800 690200 529800 691400
rect 531800 690200 532800 691400
rect 535600 689800 544200 691800
rect 545600 689800 554200 691800
rect 7200 687200 9000 688600
rect 11000 687200 12800 688600
rect 15800 687200 16800 688400
rect 18800 687200 19800 688400
rect 21800 687200 22800 688400
rect 24800 687200 25800 688400
rect 27800 687200 28800 688400
rect 30800 687200 31800 688400
rect 33800 687200 34800 688400
rect 36800 687200 37800 688400
rect 39800 687200 40800 688400
rect 42800 687200 43800 688400
rect 45800 687200 46800 688400
rect 48800 687200 49800 688400
rect 51800 687200 52800 688400
rect 54800 687200 55800 688400
rect 57800 687200 58800 688400
rect 60800 687200 61800 688400
rect 63800 687200 64800 688400
rect 66800 687200 67800 688400
rect 69800 687200 70800 688400
rect 72800 687200 73800 688400
rect 75800 687200 76800 688400
rect 78800 687200 79800 688400
rect 81800 687200 82800 688400
rect 84800 687200 85800 688400
rect 87800 687200 88800 688400
rect 90800 687200 91800 688400
rect 93800 687200 94800 688400
rect 96800 687200 97800 688400
rect 99800 687200 100800 688400
rect 102800 687200 103800 688400
rect 105800 687200 106800 688400
rect 108800 687200 109800 688400
rect 111800 687200 112800 688400
rect 114800 687200 115800 688400
rect 117800 687200 118800 688400
rect 120800 687200 121800 688400
rect 123800 687200 124800 688400
rect 126800 687200 127800 688400
rect 129800 687200 130800 688400
rect 132800 687200 133800 688400
rect 135800 687200 136800 688400
rect 138800 687200 139800 688400
rect 141800 687200 142800 688400
rect 144800 687200 145800 688400
rect 147800 687200 148800 688400
rect 150800 687200 151800 688400
rect 153800 687200 154800 688400
rect 156800 687200 157800 688400
rect 159800 687200 160800 688400
rect 162800 687200 163800 688400
rect 165800 687200 166800 688400
rect 168800 687200 169800 688400
rect 171800 687200 172800 688400
rect 174800 687200 175800 688400
rect 177800 687200 178800 688400
rect 180800 687200 181800 688400
rect 183800 687200 184800 688400
rect 186800 687200 187800 688400
rect 189800 687200 190800 688400
rect 192800 687200 193800 688400
rect 195800 687200 196800 688400
rect 198800 687200 199800 688400
rect 201800 687200 202800 688400
rect 204800 687200 205800 688400
rect 207800 687200 208800 688400
rect 210800 687200 211800 688400
rect 213800 687200 214800 688400
rect 216800 687200 217800 688400
rect 219800 687200 220800 688400
rect 222800 687200 223800 688400
rect 225800 687200 226800 688400
rect 228800 687200 229800 688400
rect 231800 687200 232800 688400
rect 234800 687200 235800 688400
rect 237800 687200 238800 688400
rect 240800 687200 241800 688400
rect 243800 687200 244800 688400
rect 246800 687200 247800 688400
rect 249800 687200 250800 688400
rect 252800 687200 253800 688400
rect 255800 687200 256800 688400
rect 258800 687200 259800 688400
rect 261800 687200 262800 688400
rect 264800 687200 265800 688400
rect 267800 687200 268800 688400
rect 270800 687200 271800 688400
rect 273800 687200 274800 688400
rect 276800 687200 277800 688400
rect 279800 687200 280800 688400
rect 282800 687200 283800 688400
rect 285800 687200 286800 688400
rect 288800 687200 289800 688400
rect 291800 687200 292800 688400
rect 294800 687200 295800 688400
rect 297800 687200 298800 688400
rect 300800 687200 301800 688400
rect 303800 687200 304800 688400
rect 306800 687200 307800 688400
rect 309800 687200 310800 688400
rect 312800 687200 313800 688400
rect 315800 687200 316800 688400
rect 318800 687200 319800 688400
rect 321800 687200 322800 688400
rect 324800 687200 325800 688400
rect 327800 687200 328800 688400
rect 330800 687200 331800 688400
rect 333800 687200 334800 688400
rect 336800 687200 337800 688400
rect 339800 687200 340800 688400
rect 342800 687200 343800 688400
rect 345800 687200 346800 688400
rect 348800 687200 349800 688400
rect 351800 687200 352800 688400
rect 354800 687200 355800 688400
rect 357800 687200 358800 688400
rect 360800 687200 361800 688400
rect 363800 687200 364800 688400
rect 366800 687200 367800 688400
rect 369800 687200 370800 688400
rect 372800 687200 373800 688400
rect 375800 687200 376800 688400
rect 378800 687200 379800 688400
rect 381800 687200 382800 688400
rect 384800 687200 385800 688400
rect 387800 687200 388800 688400
rect 390800 687200 391800 688400
rect 393800 687200 394800 688400
rect 396800 687200 397800 688400
rect 399800 687200 400800 688400
rect 402800 687200 403800 688400
rect 405800 687200 406800 688400
rect 408800 687200 409800 688400
rect 411800 687200 412800 688400
rect 414800 687200 415800 688400
rect 417800 687200 418800 688400
rect 420800 687200 421800 688400
rect 423800 687200 424800 688400
rect 426800 687200 427800 688400
rect 429800 687200 430800 688400
rect 432800 687200 433800 688400
rect 435800 687200 436800 688400
rect 438800 687200 439800 688400
rect 441800 687200 442800 688400
rect 444800 687200 445800 688400
rect 447800 687200 448800 688400
rect 450800 687200 451800 688400
rect 453800 687200 454800 688400
rect 456800 687200 457800 688400
rect 459800 687200 460800 688400
rect 462800 687200 463800 688400
rect 465800 687200 466800 688400
rect 468800 687200 469800 688400
rect 471800 687200 472800 688400
rect 474800 687200 475800 688400
rect 477800 687200 478800 688400
rect 480800 687200 481800 688400
rect 483800 687200 484800 688400
rect 486800 687200 487800 688400
rect 489800 687200 490800 688400
rect 492800 687200 493800 688400
rect 495800 687200 496800 688400
rect 498800 687200 499800 688400
rect 501800 687200 502800 688400
rect 504800 687200 505800 688400
rect 507800 687200 508800 688400
rect 510800 687200 511800 688400
rect 513800 687200 514800 688400
rect 516800 687200 517800 688400
rect 519800 687200 520800 688400
rect 522800 687200 523800 688400
rect 525800 687200 526800 688400
rect 528800 687200 529800 688400
rect 531800 687200 532800 688400
rect 535600 685800 544200 687800
rect 545600 685800 554200 687800
rect 7200 684200 9000 685600
rect 11000 684200 12800 685600
rect 15800 684200 16800 685400
rect 18800 684200 19800 685400
rect 21800 684200 22800 685400
rect 24800 684200 25800 685400
rect 27800 684200 28800 685400
rect 30800 684200 31800 685400
rect 33800 684200 34800 685400
rect 36800 684200 37800 685400
rect 39800 684200 40800 685400
rect 42800 684200 43800 685400
rect 45800 684200 46800 685400
rect 48800 684200 49800 685400
rect 51800 684200 52800 685400
rect 54800 684200 55800 685400
rect 57800 684200 58800 685400
rect 60800 684200 61800 685400
rect 63800 684200 64800 685400
rect 66800 684200 67800 685400
rect 69800 684200 70800 685400
rect 72800 684200 73800 685400
rect 75800 684200 76800 685400
rect 78800 684200 79800 685400
rect 81800 684200 82800 685400
rect 84800 684200 85800 685400
rect 87800 684200 88800 685400
rect 90800 684200 91800 685400
rect 93800 684200 94800 685400
rect 96800 684200 97800 685400
rect 99800 684200 100800 685400
rect 102800 684200 103800 685400
rect 105800 684200 106800 685400
rect 108800 684200 109800 685400
rect 111800 684200 112800 685400
rect 114800 684200 115800 685400
rect 117800 684200 118800 685400
rect 120800 684200 121800 685400
rect 123800 684200 124800 685400
rect 126800 684200 127800 685400
rect 129800 684200 130800 685400
rect 132800 684200 133800 685400
rect 135800 684200 136800 685400
rect 138800 684200 139800 685400
rect 141800 684200 142800 685400
rect 144800 684200 145800 685400
rect 147800 684200 148800 685400
rect 150800 684200 151800 685400
rect 153800 684200 154800 685400
rect 156800 684200 157800 685400
rect 159800 684200 160800 685400
rect 162800 684200 163800 685400
rect 165800 684200 166800 685400
rect 168800 684200 169800 685400
rect 171800 684200 172800 685400
rect 174800 684200 175800 685400
rect 177800 684200 178800 685400
rect 180800 684200 181800 685400
rect 183800 684200 184800 685400
rect 186800 684200 187800 685400
rect 189800 684200 190800 685400
rect 192800 684200 193800 685400
rect 195800 684200 196800 685400
rect 198800 684200 199800 685400
rect 201800 684200 202800 685400
rect 204800 684200 205800 685400
rect 207800 684200 208800 685400
rect 210800 684200 211800 685400
rect 213800 684200 214800 685400
rect 216800 684200 217800 685400
rect 219800 684200 220800 685400
rect 222800 684200 223800 685400
rect 225800 684200 226800 685400
rect 228800 684200 229800 685400
rect 231800 684200 232800 685400
rect 234800 684200 235800 685400
rect 237800 684200 238800 685400
rect 240800 684200 241800 685400
rect 243800 684200 244800 685400
rect 246800 684200 247800 685400
rect 249800 684200 250800 685400
rect 252800 684200 253800 685400
rect 255800 684200 256800 685400
rect 258800 684200 259800 685400
rect 261800 684200 262800 685400
rect 264800 684200 265800 685400
rect 267800 684200 268800 685400
rect 270800 684200 271800 685400
rect 273800 684200 274800 685400
rect 276800 684200 277800 685400
rect 279800 684200 280800 685400
rect 282800 684200 283800 685400
rect 285800 684200 286800 685400
rect 288800 684200 289800 685400
rect 291800 684200 292800 685400
rect 294800 684200 295800 685400
rect 297800 684200 298800 685400
rect 300800 684200 301800 685400
rect 303800 684200 304800 685400
rect 306800 684200 307800 685400
rect 309800 684200 310800 685400
rect 312800 684200 313800 685400
rect 315800 684200 316800 685400
rect 318800 684200 319800 685400
rect 321800 684200 322800 685400
rect 324800 684200 325800 685400
rect 327800 684200 328800 685400
rect 330800 684200 331800 685400
rect 333800 684200 334800 685400
rect 336800 684200 337800 685400
rect 339800 684200 340800 685400
rect 342800 684200 343800 685400
rect 345800 684200 346800 685400
rect 348800 684200 349800 685400
rect 351800 684200 352800 685400
rect 354800 684200 355800 685400
rect 357800 684200 358800 685400
rect 360800 684200 361800 685400
rect 363800 684200 364800 685400
rect 366800 684200 367800 685400
rect 369800 684200 370800 685400
rect 372800 684200 373800 685400
rect 375800 684200 376800 685400
rect 378800 684200 379800 685400
rect 381800 684200 382800 685400
rect 384800 684200 385800 685400
rect 387800 684200 388800 685400
rect 390800 684200 391800 685400
rect 393800 684200 394800 685400
rect 396800 684200 397800 685400
rect 399800 684200 400800 685400
rect 402800 684200 403800 685400
rect 405800 684200 406800 685400
rect 408800 684200 409800 685400
rect 411800 684200 412800 685400
rect 414800 684200 415800 685400
rect 417800 684200 418800 685400
rect 420800 684200 421800 685400
rect 423800 684200 424800 685400
rect 426800 684200 427800 685400
rect 429800 684200 430800 685400
rect 432800 684200 433800 685400
rect 435800 684200 436800 685400
rect 438800 684200 439800 685400
rect 441800 684200 442800 685400
rect 444800 684200 445800 685400
rect 447800 684200 448800 685400
rect 450800 684200 451800 685400
rect 453800 684200 454800 685400
rect 456800 684200 457800 685400
rect 459800 684200 460800 685400
rect 462800 684200 463800 685400
rect 465800 684200 466800 685400
rect 468800 684200 469800 685400
rect 471800 684200 472800 685400
rect 474800 684200 475800 685400
rect 477800 684200 478800 685400
rect 480800 684200 481800 685400
rect 483800 684200 484800 685400
rect 486800 684200 487800 685400
rect 489800 684200 490800 685400
rect 492800 684200 493800 685400
rect 495800 684200 496800 685400
rect 498800 684200 499800 685400
rect 501800 684200 502800 685400
rect 504800 684200 505800 685400
rect 507800 684200 508800 685400
rect 510800 684200 511800 685400
rect 513800 684200 514800 685400
rect 516800 684200 517800 685400
rect 519800 684200 520800 685400
rect 522800 684200 523800 685400
rect 525800 684200 526800 685400
rect 528800 684200 529800 685400
rect 531800 684200 532800 685400
rect 7200 681200 9000 682600
rect 11000 681200 12800 682600
rect 15800 681200 16800 682400
rect 18800 681200 19800 682400
rect 21800 681200 22800 682400
rect 24800 681200 25800 682400
rect 27800 681200 28800 682400
rect 30800 681200 31800 682400
rect 33800 681200 34800 682400
rect 36800 681200 37800 682400
rect 39800 681200 40800 682400
rect 42800 681200 43800 682400
rect 45800 681200 46800 682400
rect 48800 681200 49800 682400
rect 51800 681200 52800 682400
rect 54800 681200 55800 682400
rect 57800 681200 58800 682400
rect 60800 681200 61800 682400
rect 63800 681200 64800 682400
rect 66800 681200 67800 682400
rect 69800 681200 70800 682400
rect 72800 681200 73800 682400
rect 75800 681200 76800 682400
rect 78800 681200 79800 682400
rect 81800 681200 82800 682400
rect 84800 681200 85800 682400
rect 87800 681200 88800 682400
rect 90800 681200 91800 682400
rect 93800 681200 94800 682400
rect 96800 681200 97800 682400
rect 99800 681200 100800 682400
rect 102800 681200 103800 682400
rect 105800 681200 106800 682400
rect 108800 681200 109800 682400
rect 111800 681200 112800 682400
rect 114800 681200 115800 682400
rect 117800 681200 118800 682400
rect 120800 681200 121800 682400
rect 123800 681200 124800 682400
rect 126800 681200 127800 682400
rect 129800 681200 130800 682400
rect 132800 681200 133800 682400
rect 135800 681200 136800 682400
rect 138800 681200 139800 682400
rect 141800 681200 142800 682400
rect 144800 681200 145800 682400
rect 147800 681200 148800 682400
rect 150800 681200 151800 682400
rect 153800 681200 154800 682400
rect 156800 681200 157800 682400
rect 159800 681200 160800 682400
rect 162800 681200 163800 682400
rect 165800 681200 166800 682400
rect 168800 681200 169800 682400
rect 171800 681200 172800 682400
rect 174800 681200 175800 682400
rect 177800 681200 178800 682400
rect 180800 681200 181800 682400
rect 183800 681200 184800 682400
rect 186800 681200 187800 682400
rect 189800 681200 190800 682400
rect 192800 681200 193800 682400
rect 195800 681200 196800 682400
rect 198800 681200 199800 682400
rect 201800 681200 202800 682400
rect 204800 681200 205800 682400
rect 207800 681200 208800 682400
rect 210800 681200 211800 682400
rect 213800 681200 214800 682400
rect 216800 681200 217800 682400
rect 219800 681200 220800 682400
rect 222800 681200 223800 682400
rect 225800 681200 226800 682400
rect 228800 681200 229800 682400
rect 231800 681200 232800 682400
rect 234800 681200 235800 682400
rect 237800 681200 238800 682400
rect 240800 681200 241800 682400
rect 243800 681200 244800 682400
rect 246800 681200 247800 682400
rect 249800 681200 250800 682400
rect 252800 681200 253800 682400
rect 255800 681200 256800 682400
rect 258800 681200 259800 682400
rect 261800 681200 262800 682400
rect 264800 681200 265800 682400
rect 267800 681200 268800 682400
rect 270800 681200 271800 682400
rect 273800 681200 274800 682400
rect 276800 681200 277800 682400
rect 279800 681200 280800 682400
rect 282800 681200 283800 682400
rect 285800 681200 286800 682400
rect 288800 681200 289800 682400
rect 291800 681200 292800 682400
rect 294800 681200 295800 682400
rect 297800 681200 298800 682400
rect 300800 681200 301800 682400
rect 303800 681200 304800 682400
rect 306800 681200 307800 682400
rect 309800 681200 310800 682400
rect 312800 681200 313800 682400
rect 315800 681200 316800 682400
rect 318800 681200 319800 682400
rect 321800 681200 322800 682400
rect 324800 681200 325800 682400
rect 327800 681200 328800 682400
rect 330800 681200 331800 682400
rect 333800 681200 334800 682400
rect 336800 681200 337800 682400
rect 339800 681200 340800 682400
rect 342800 681200 343800 682400
rect 345800 681200 346800 682400
rect 348800 681200 349800 682400
rect 351800 681200 352800 682400
rect 354800 681200 355800 682400
rect 357800 681200 358800 682400
rect 360800 681200 361800 682400
rect 363800 681200 364800 682400
rect 366800 681200 367800 682400
rect 369800 681200 370800 682400
rect 372800 681200 373800 682400
rect 375800 681200 376800 682400
rect 378800 681200 379800 682400
rect 381800 681200 382800 682400
rect 384800 681200 385800 682400
rect 387800 681200 388800 682400
rect 390800 681200 391800 682400
rect 393800 681200 394800 682400
rect 396800 681200 397800 682400
rect 399800 681200 400800 682400
rect 402800 681200 403800 682400
rect 405800 681200 406800 682400
rect 408800 681200 409800 682400
rect 411800 681200 412800 682400
rect 414800 681200 415800 682400
rect 417800 681200 418800 682400
rect 420800 681200 421800 682400
rect 423800 681200 424800 682400
rect 426800 681200 427800 682400
rect 429800 681200 430800 682400
rect 432800 681200 433800 682400
rect 435800 681200 436800 682400
rect 438800 681200 439800 682400
rect 441800 681200 442800 682400
rect 444800 681200 445800 682400
rect 447800 681200 448800 682400
rect 450800 681200 451800 682400
rect 453800 681200 454800 682400
rect 456800 681200 457800 682400
rect 459800 681200 460800 682400
rect 462800 681200 463800 682400
rect 465800 681200 466800 682400
rect 468800 681200 469800 682400
rect 471800 681200 472800 682400
rect 474800 681200 475800 682400
rect 477800 681200 478800 682400
rect 480800 681200 481800 682400
rect 483800 681200 484800 682400
rect 486800 681200 487800 682400
rect 489800 681200 490800 682400
rect 492800 681200 493800 682400
rect 495800 681200 496800 682400
rect 498800 681200 499800 682400
rect 501800 681200 502800 682400
rect 504800 681200 505800 682400
rect 507800 681200 508800 682400
rect 510800 681200 511800 682400
rect 513800 681200 514800 682400
rect 516800 681200 517800 682400
rect 519800 681200 520800 682400
rect 522800 681200 523800 682400
rect 525800 681200 526800 682400
rect 528800 681200 529800 682400
rect 531800 681200 532800 682400
rect 535600 681800 544200 683800
rect 545600 681800 554200 683800
rect 7200 678200 9000 679600
rect 11000 678200 12800 679600
rect 7200 675200 9000 676600
rect 11000 675200 12800 676600
rect 7200 672200 9000 673600
rect 11000 672200 12800 673600
rect 7200 669200 9000 670600
rect 11000 669200 12800 670600
rect 7200 666200 9000 667600
rect 11000 666200 12800 667600
rect 7200 663200 9000 664600
rect 11000 663200 12800 664600
rect 7200 660200 9000 661600
rect 11000 660200 12800 661600
rect 7200 657200 9000 658600
rect 11000 657200 12800 658600
rect 4800 654800 6200 656000
rect 7200 654200 9000 655600
rect 11000 654200 12800 655600
rect 4800 652800 6200 654000
rect 4800 650800 6200 652000
rect 7200 651200 9000 652600
rect 11000 651200 12800 652600
rect 4800 648800 6200 650000
rect 7200 648200 9000 649600
rect 11000 648200 12800 649600
rect 4800 646800 6200 648000
rect 4800 644800 6200 646000
rect 7200 645200 9000 646600
rect 11000 645200 12800 646600
rect 4800 642800 6200 644000
rect 7200 642200 9000 643600
rect 11000 642200 12800 643600
rect 4800 640800 6200 642000
rect 4800 638800 6200 640000
rect 7200 639200 9000 640600
rect 11000 639200 12800 640600
rect 4800 636800 6200 638000
rect 7200 636200 9000 637600
rect 11000 636200 12800 637600
rect 4800 634800 6200 636000
rect 4800 632800 6200 634000
rect 7200 633200 9000 634600
rect 11000 633200 12800 634600
rect 4800 630800 6200 632000
rect 7400 630800 8800 632000
rect 475800 676000 477200 677400
rect 535600 677800 544200 679800
rect 545600 677800 554200 679800
rect 475800 674000 477200 675400
rect 475800 672000 477200 673400
rect 475800 670000 477200 671400
rect 475800 668000 477200 669400
rect 475800 666000 477200 667400
rect 475800 664000 477200 665400
rect 475800 662000 477200 663400
rect 475800 660000 477200 661400
rect 475800 658000 477200 659400
rect 475800 656000 477200 657400
rect 475800 654000 477200 655400
rect 475800 652000 477200 653400
rect 475800 650000 477200 651400
rect 475800 648000 477200 649400
rect 475800 646000 477200 647400
rect 475800 644000 477200 645400
rect 535600 673800 544200 675800
rect 545600 673800 554200 675800
rect 520580 664340 526480 669740
rect 535600 669800 544200 671800
rect 545600 669800 554200 671800
rect 535600 665800 544200 667800
rect 545600 665800 554200 667800
rect 535600 661800 544200 663800
rect 545600 661800 554200 663800
rect 475800 642000 477200 643400
rect 475800 640000 477200 641400
rect 475800 638000 477200 639400
rect 475800 636000 477200 637400
rect 475800 634000 477200 635400
rect 475800 632000 477200 633400
rect 4800 628800 6200 630000
rect 7400 628800 8800 630000
rect 4800 626800 6200 628000
rect 7400 626800 8800 628000
rect 4800 624800 6200 626000
rect 7400 624800 8800 626000
rect 4800 622800 6200 624000
rect 7400 622800 8800 624000
rect 4800 620800 6200 622000
rect 7400 620800 8800 622000
rect 4800 618800 6200 620000
rect 7400 618800 8800 620000
rect 4800 616800 6200 618000
rect 7400 616800 8800 618000
rect 4800 614800 6200 616000
rect 7400 614800 8800 616000
rect 4800 612800 6200 614000
rect 7400 612800 8800 614000
rect 4800 610800 6200 612000
rect 7400 610800 8800 612000
rect 4800 608800 6200 610000
rect 7400 608800 8800 610000
rect 4800 606800 6200 608000
rect 7400 606800 8800 608000
rect 4800 604800 6200 606000
rect 7400 604800 8800 606000
rect 4800 602800 6200 604000
rect 7400 602800 8800 604000
rect 4800 600800 6200 602000
rect 7400 600800 8800 602000
rect 4800 598800 6200 600000
rect 7400 598800 8800 600000
rect 4800 596800 6200 598000
rect 7400 596800 8800 598000
rect 4800 594800 6200 596000
rect 7400 594800 8800 596000
rect 4800 592800 6200 594000
rect 7400 592800 8800 594000
rect 4800 590800 6200 592000
rect 7400 590800 8800 592000
rect 4800 588800 6200 590000
rect 7400 588800 8800 590000
rect 4800 586800 6200 588000
rect 7400 586800 8800 588000
rect 4800 584800 6200 586000
rect 7400 584800 8800 586000
rect 4800 582800 6200 584000
rect 7400 582800 8800 584000
rect 4800 580800 6200 582000
rect 7400 580800 8800 582000
rect 4800 578800 6200 580000
rect 7400 578800 8800 580000
rect 4800 576800 6200 578000
rect 7400 576800 8800 578000
rect 4800 574800 6200 576000
rect 7400 574800 8800 576000
rect 4800 572800 6200 574000
rect 7400 572800 8800 574000
rect 4800 570800 6200 572000
rect 7400 570800 8800 572000
rect 4800 568800 6200 570000
rect 7400 568800 8800 570000
rect 4800 566800 6200 568000
rect 7400 566800 8800 568000
rect 4800 564800 6200 566000
rect 7400 564800 8800 566000
rect 870 549250 2600 564320
rect 16000 629600 16800 630200
rect 16000 626600 16800 627200
rect 16000 623600 16800 624200
rect 16000 620600 16800 621200
rect 16000 617600 16800 618200
rect 16000 614600 16800 615200
rect 16000 611600 16800 612200
rect 16000 608600 16800 609200
rect 16000 605600 16800 606200
rect 16000 602600 16800 603200
rect 16000 599600 16800 600200
rect 16000 596600 16800 597200
rect 16000 593600 16800 594200
rect 16000 590600 16800 591200
rect 16000 587600 16800 588200
rect 16000 584600 16800 585200
rect 16000 581600 16800 582200
rect 16000 578600 16800 579200
rect 16000 575600 16800 576200
rect 16000 572600 16800 573200
rect 16000 569600 16800 570200
rect 16000 566600 16800 567200
rect 475800 630000 477200 631400
rect 475800 628000 477200 629400
rect 475800 626000 477200 627400
rect 535600 657800 544200 659800
rect 545600 657800 554200 659800
rect 535600 653800 544200 655800
rect 545600 653800 554200 655800
rect 535600 649800 544200 651800
rect 545600 649800 554200 651800
rect 520780 641340 526680 646740
rect 535600 645800 544200 647800
rect 545600 645800 554200 647800
rect 535600 641800 544200 643800
rect 545600 641800 554200 643800
rect 535600 637800 544200 639800
rect 545600 637800 554200 639800
rect 535600 633800 544200 635800
rect 545600 633800 554200 635800
rect 499340 628360 507010 629510
rect 535600 629800 544200 631800
rect 545600 629800 554200 631800
rect 576690 630020 583530 644270
rect 475800 624000 477200 625400
rect 475800 622000 477200 623400
rect 475800 620000 477200 621400
rect 475800 618000 477200 619400
rect 475800 616000 477200 617400
rect 520580 617740 526580 623040
rect 475800 614000 477200 615400
rect 475800 612000 477200 613400
rect 475800 610000 477200 611400
rect 475800 608000 477200 609400
rect 475800 606000 477200 607400
rect 475800 604000 477200 605400
rect 475800 602000 477200 603400
rect 475800 600000 477200 601400
rect 475800 598000 477200 599400
rect 475800 596000 477200 597400
rect 475800 594000 477200 595400
rect 475800 592000 477200 593400
rect 475800 590000 477200 591400
rect 475800 588000 477200 589400
rect 475800 586000 477200 587400
rect 475800 584000 477200 585400
rect 475800 582000 477200 583400
rect 475800 580000 477200 581400
rect 475800 578000 477200 579400
rect 475800 576000 477200 577400
rect 475800 574000 477200 575400
rect 475800 572000 477200 573400
rect 475800 570000 477200 571400
rect 475800 568000 477200 569400
rect 475800 566000 477200 567400
rect 4800 562800 6200 564000
rect 7400 562800 8800 564000
rect 4800 560800 6200 562000
rect 7400 560800 8800 562000
rect 4800 558800 6200 560000
rect 7400 558800 8800 560000
rect 4800 556800 6200 558000
rect 7400 556800 8800 558000
rect 4800 554800 6200 556000
rect 7400 554800 8800 556000
rect 4800 552800 6200 554000
rect 7400 552800 8800 554000
rect 4800 550800 6200 552000
rect 7400 550800 8800 552000
rect 4800 548800 6200 550000
rect 7400 548800 8800 550000
rect 4800 546800 6200 548000
rect 7400 546800 8800 548000
rect 4800 544800 6200 546000
rect 7400 544800 8800 546000
rect 4800 542800 6200 544000
rect 7400 542800 8800 544000
rect 4800 540800 6200 542000
rect 7400 540800 8800 542000
rect 4800 538800 6200 540000
rect 7400 538800 8800 540000
rect 16000 563600 16800 564200
rect 16000 560600 16800 561200
rect 16000 558000 16800 558200
rect 16000 557600 16800 558000
rect 16000 554800 16800 555200
rect 16000 554600 16800 554800
rect 16000 551600 16800 552200
rect 16000 548800 16800 549200
rect 16000 548600 16800 548800
rect 16000 547200 16800 547800
rect 16000 544200 16800 544800
rect 475800 564000 477200 565400
rect 475800 562000 477200 563400
rect 475800 560000 477200 561400
rect 512590 568680 518490 574080
rect 475800 558000 477200 559400
rect 475800 556000 477200 557400
rect 475800 554000 477200 555400
rect 475800 552000 477200 553400
rect 475800 550000 477200 551400
rect 475800 548000 477200 549400
rect 475800 546000 477200 547400
rect 475800 544000 477200 545400
rect 16000 541200 16800 541800
rect 16000 538200 16800 538800
rect 3800 536400 5200 537600
rect 3800 534400 5200 535600
rect 16000 535200 16800 535800
rect 3800 532400 5200 533600
rect 3800 531120 5200 531600
rect 3800 530740 4130 531120
rect 4130 530740 4920 531120
rect 4920 530740 5200 531120
rect 3800 530400 5200 530740
rect 3800 529050 5200 529600
rect 3800 528670 4130 529050
rect 4130 528670 4920 529050
rect 4920 528670 5200 529050
rect 3800 528400 5200 528670
rect 3800 526400 5200 527600
rect 15800 531800 17100 532200
rect 15800 531100 17100 531500
rect 15800 530500 17100 530900
rect 15800 529800 17100 530200
rect 15800 529100 17100 529500
rect 15800 528400 17100 528800
rect 3800 524400 5200 525600
rect 3800 522400 5200 523600
rect 3800 520400 5200 521600
rect 3800 518400 5200 519600
rect 3800 516400 5200 517600
rect 3800 514400 5200 515600
rect 3800 512400 5200 513600
rect 3800 510400 5200 511600
rect 3800 508400 5200 509600
rect 3800 506400 5200 507600
rect 3800 504400 5200 505600
rect 3800 502400 5200 503600
rect 3800 500400 5200 501600
rect 3800 498400 5200 499600
rect 3800 496400 5200 497600
rect 3800 494400 5200 495600
rect 3800 492400 5200 493600
rect 3800 490400 5200 491600
rect 3800 488400 5200 489600
rect 3800 486400 5200 487600
rect 3800 484400 5200 485600
rect 3800 482400 5200 483600
rect 3800 480400 5200 481600
rect 3800 478400 5200 479600
rect 3800 476400 5200 477600
rect 3800 474400 5200 475600
rect 3800 472400 5200 473600
rect 3800 470400 5200 471600
rect 3800 468400 5200 469600
rect 3800 466400 5200 467600
rect 3800 464400 5200 465600
rect 3800 462400 5200 463600
rect 3800 460400 5200 461600
rect 3800 458400 5200 459600
rect 3800 456400 5200 457600
rect 3800 454400 5200 455600
rect 3800 452400 5200 453600
rect 3800 450400 5200 451600
rect 3800 448400 5200 449600
rect 3800 446400 5200 447600
rect 3800 444400 5200 445600
rect 3800 442400 5200 443600
rect 3800 440400 5200 441600
rect 3800 438400 5200 439600
rect 3800 436400 5200 437600
rect 3800 434400 5200 435600
rect 3800 432400 5200 433600
rect 16000 526600 16800 527200
rect 16000 523600 16800 524200
rect 16000 520600 16800 521200
rect 16000 517600 16800 518200
rect 16000 514600 16800 515200
rect 16000 511600 16800 512200
rect 16000 508600 16800 509200
rect 16000 505600 16800 506200
rect 16000 502600 16800 503200
rect 16000 499600 16800 500200
rect 16000 496600 16800 497200
rect 16000 493600 16800 494200
rect 16000 490600 16800 491200
rect 16000 487600 16800 488200
rect 16000 484600 16800 485200
rect 16000 481600 16800 482200
rect 16000 478600 16800 479200
rect 16000 475600 16800 476200
rect 16000 472600 16800 473200
rect 16000 469600 16800 470200
rect 16000 466600 16800 467200
rect 16000 463600 16800 464200
rect 16000 460600 16800 461200
rect 16000 457600 16800 458200
rect 16000 454600 16800 455200
rect 16000 451600 16800 452200
rect 16000 448600 16800 449200
rect 16000 445600 16800 446200
rect 16000 442600 16800 443200
rect 16000 439600 16800 440200
rect 16000 436600 16800 437200
rect 16000 433600 16800 434200
rect 16000 430600 16800 431200
rect 16000 427600 16800 428200
rect 16000 424600 16800 425200
rect 16000 421600 16800 422200
rect 16000 418600 16800 419200
rect 16000 415600 16800 416200
rect 16000 412600 16800 413200
rect 16000 409600 16800 410200
rect 16000 406600 16800 407200
rect 16000 403600 16800 404200
rect 16000 400600 16800 401200
rect 16000 397600 16800 398200
rect 16000 394600 16800 395200
rect 16000 391600 16800 392200
rect 16000 388600 16800 389200
rect 16000 385600 16800 386200
rect 16000 382600 16800 383200
rect 16000 379600 16800 380200
rect 16000 376600 16800 377200
rect 1000 375000 2000 375400
rect 1000 374400 2000 374800
rect 1000 373600 2000 374000
rect 1000 372800 2000 373200
rect 1000 372000 2000 372400
rect 1000 371200 2000 371600
rect 1000 370400 2000 370800
rect 16000 373600 16800 374200
rect 16000 370600 16800 371200
rect 800 368800 1400 369400
rect 800 366800 1400 367400
rect 800 364800 1400 365400
rect 800 362800 1400 363400
rect 800 360800 1400 361400
rect 800 358800 1400 359400
rect 800 356800 1400 357400
rect 800 354800 1400 355400
rect 800 352800 1400 353400
rect 800 350800 1400 351400
rect 800 348800 1400 349400
rect 800 346800 1400 347400
rect 800 344800 1400 345400
rect 16000 341200 16800 341800
rect 16000 338200 16800 338800
rect 16000 335200 16800 335800
rect 16000 332200 16800 332800
rect 475800 542000 477200 543400
rect 475800 540000 477200 541400
rect 475800 538000 477200 539400
rect 475800 536000 477200 537400
rect 475800 534000 477200 535400
rect 565180 568810 571080 574210
rect 512790 545680 518690 551080
rect 475800 532000 477200 533400
rect 491350 532700 499020 533850
rect 565380 545810 571280 551210
rect 475800 530000 477200 531400
rect 475800 528000 477200 529400
rect 475800 526000 477200 527400
rect 475800 524000 477200 525400
rect 475800 522000 477200 523400
rect 475800 520000 477200 521400
rect 512590 522080 518590 527380
rect 475800 518000 477200 519400
rect 475800 516000 477200 517400
rect 543940 532830 551610 533980
rect 565180 522210 571180 527510
rect 475800 514000 477200 515400
rect 475800 512000 477200 513400
rect 475800 510000 477200 511400
rect 475800 508000 477200 509400
rect 475800 506000 477200 507400
rect 475800 504000 477200 505400
rect 475800 502000 477200 503400
rect 475800 500000 477200 501400
rect 475800 498000 477200 499400
rect 475800 496000 477200 497400
rect 475800 494000 477200 495400
rect 475800 492000 477200 493400
rect 529410 493080 530560 500750
rect 475800 490000 477200 491400
rect 475800 488000 477200 489400
rect 475800 486000 477200 487400
rect 475800 484000 477200 485400
rect 475800 482000 477200 483400
rect 475800 480000 477200 481400
rect 475800 478000 477200 479400
rect 475800 476000 477200 477400
rect 475800 474000 477200 475400
rect 475800 472000 477200 473400
rect 518790 473510 524090 479510
rect 542390 473410 547790 479310
rect 565390 473610 570790 479510
rect 475800 470000 477200 471400
rect 475800 468000 477200 469400
rect 475800 466000 477200 467400
rect 475800 464000 477200 465400
rect 475800 462000 477200 463400
rect 475800 460000 477200 461400
rect 475800 458000 477200 459400
rect 475800 456000 477200 457400
rect 475800 454000 477200 455400
rect 475800 452000 477200 453400
rect 475800 450000 477200 451400
rect 475800 448000 477200 449400
rect 475800 446000 477200 447400
rect 475800 444000 477200 445400
rect 475800 442000 477200 443400
rect 475800 440000 477200 441400
rect 475800 438000 477200 439400
rect 475800 436000 477200 437400
rect 475800 434000 477200 435400
rect 475800 432000 477200 433400
rect 475800 430000 477200 431400
rect 475800 428000 477200 429400
rect 475800 426000 477200 427400
rect 475800 424000 477200 425400
rect 475800 422000 477200 423400
rect 475800 420000 477200 421400
rect 475800 418000 477200 419400
rect 475800 416000 477200 417400
rect 475800 414000 477200 415400
rect 475800 412000 477200 413400
rect 475800 410000 477200 411400
rect 475800 408000 477200 409400
rect 475800 406000 477200 407400
rect 475800 404000 477200 405400
rect 475800 402000 477200 403400
rect 475800 400000 477200 401400
rect 475800 398000 477200 399400
rect 475800 396000 477200 397400
rect 475800 394000 477200 395400
rect 475800 392000 477200 393400
rect 475800 390000 477200 391400
rect 475800 388000 477200 389400
rect 475800 386000 477200 387400
rect 475800 384000 477200 385400
rect 475800 382000 477200 383400
rect 475800 380000 477200 381400
rect 475800 378000 477200 379400
rect 475800 376000 477200 377400
rect 475800 374000 477200 375400
rect 475800 372000 477200 373400
rect 475800 370000 477200 371400
rect 475800 368000 477200 369400
rect 475800 366000 477200 367400
rect 475800 364000 477200 365400
rect 475800 362000 477200 363400
rect 475800 360000 477200 361400
rect 475800 358000 477200 359400
rect 475800 356000 477200 357400
rect 475800 354000 477200 355400
rect 475800 352000 477200 353400
rect 475800 350000 477200 351400
rect 475800 348000 477200 349400
rect 475800 346000 477200 347400
rect 475800 344000 477200 345400
rect 475800 342000 477200 343400
rect 475800 340000 477200 341400
rect 475800 338000 477200 339400
rect 475800 336000 477200 337400
rect 475800 334000 477200 335400
rect 475800 332000 477200 333400
rect 16000 329200 16800 329800
rect 16000 326200 16800 326800
rect 16000 323200 16800 323800
rect 16000 320200 16800 320800
rect 16000 317200 16800 317800
rect 16000 314200 16800 314800
rect 16000 311200 16800 311800
rect 16000 308200 16800 308800
rect 16000 305200 16800 305800
rect 16000 302200 16800 302800
rect 16000 299200 16800 299800
rect 16000 296200 16800 296800
rect 16000 293200 16800 293800
rect 16000 290200 16800 290800
rect 16000 287200 16800 287800
rect 16000 284200 16800 284800
rect 16000 281200 16800 281800
rect 16000 278200 16800 278800
rect 16000 275200 16800 275800
rect 16000 272200 16800 272800
rect 16000 269200 16800 269800
rect 16000 266200 16800 266800
rect 16000 263200 16800 263800
rect 16000 260200 16800 260800
rect 16000 257200 16800 257800
rect 16000 254200 16800 254800
rect 16000 251200 16800 251800
rect 16000 248200 16800 248800
rect 16000 245200 16800 245800
rect 16000 242200 16800 242800
rect 16000 239200 16800 239800
rect 16000 236200 16800 236800
rect 16000 233200 16800 233800
rect 16000 230200 16800 230800
rect 16000 227200 16800 227800
rect 16000 224200 16800 224800
rect 16000 221200 16800 221800
rect 16000 218200 16800 218800
rect 16000 215200 16800 215800
rect 16000 212200 16800 212800
rect 16000 209200 16800 209800
rect 16000 206200 16800 206800
rect 16000 203200 16800 203800
rect 16000 200200 16800 200800
rect 16000 197200 16800 197800
rect 16000 194200 16800 194800
rect 16000 191200 16800 191800
rect 16000 188200 16800 188800
rect 16000 185200 16800 185800
rect 16000 182200 16800 182800
rect 16000 179200 16800 179800
rect 700 163110 2330 177370
rect 16000 176200 16800 176800
rect 16000 173200 16800 173800
rect 16000 170200 16800 170800
rect 16000 167200 16800 167800
rect 16000 164200 16800 164800
rect 16000 161200 16800 161800
rect 16000 158200 16800 158800
rect 16000 155200 16800 155800
rect 16000 152200 16800 152800
rect 16000 149200 16800 149800
rect 16000 146200 16800 146800
rect 16000 143200 16800 143800
rect 16000 140200 16800 140800
rect 16000 137200 16800 137800
rect 16000 134200 16800 134800
rect 16000 131200 16800 131800
rect 16000 128200 16800 128800
rect 16000 125200 16800 125800
rect 16000 122200 16800 122800
rect 16000 119200 16800 119800
rect 16000 116200 16800 116800
rect 16000 113200 16800 113800
rect 16000 110200 16800 110800
rect 16000 107200 16800 107800
rect 16000 104200 16800 104800
rect 16000 101200 16800 101800
rect 16000 98200 16800 98800
rect 16000 95200 16800 95800
rect 16000 92200 16800 92800
rect 16000 89200 16800 89800
rect 16000 86200 16800 86800
rect 16000 83200 16800 83800
rect 16000 80200 16800 80800
rect 16000 77200 16800 77800
rect 16000 74200 16800 74800
rect 16000 71200 16800 71800
rect 16000 68200 16800 68800
rect 16000 65200 16800 65800
rect 16000 62200 16800 62800
rect 16000 59200 16800 59800
rect 16000 56200 16800 56800
rect 16000 53200 16800 53800
rect 16000 50200 16800 50800
rect 16000 47200 16800 47800
rect 16000 44200 16800 44800
rect 16000 41200 16800 41800
rect 16000 38200 16800 38800
rect 16000 35200 16800 35800
rect 16000 32200 16800 32800
rect 16000 29200 16800 29800
rect 16000 26200 16800 26800
rect 16000 23200 16800 23800
rect 16000 20200 16800 20800
rect 16000 17200 16800 17800
rect 16000 14200 16800 14800
rect 16000 11200 16800 11800
rect 16000 8200 16800 8800
rect 16000 5200 16800 5800
rect 475800 330000 477200 331400
rect 475800 328000 477200 329400
rect 475800 326000 477200 327400
rect 475800 324000 477200 325400
rect 475800 322000 477200 323400
rect 475800 320000 477200 321400
rect 475800 318000 477200 319400
rect 475800 316000 477200 317400
rect 475800 314000 477200 315400
rect 475800 312000 477200 313400
rect 475800 310000 477200 311400
rect 475800 308000 477200 309400
rect 475800 306000 477200 307400
rect 475800 304000 477200 305400
rect 475800 302000 477200 303400
rect 475800 300000 477200 301400
rect 475800 298000 477200 299400
rect 475800 296000 477200 297400
rect 475800 294000 477200 295400
rect 475800 292000 477200 293400
rect 475800 290000 477200 291400
rect 475800 288000 477200 289400
rect 475800 286000 477200 287400
rect 475800 284000 477200 285400
rect 475800 282000 477200 283400
rect 475800 280000 477200 281400
rect 475800 278000 477200 279400
rect 475800 276000 477200 277400
rect 475800 274000 477200 275400
rect 475800 272000 477200 273400
rect 475800 270000 477200 271400
rect 475800 268000 477200 269400
rect 475800 266000 477200 267400
rect 475800 264000 477200 265400
rect 475800 262000 477200 263400
rect 475800 260000 477200 261400
rect 475800 258000 477200 259400
rect 576800 395800 582200 396400
rect 576800 393800 582200 394400
rect 576800 391800 582200 392400
rect 576800 389800 582200 390400
rect 576800 387800 582200 388400
rect 576800 385800 582200 386400
rect 576800 383800 582200 384400
rect 576800 381800 582200 382400
rect 576800 379800 582200 380400
rect 576800 377800 582200 378400
rect 576800 375800 582200 376400
rect 576800 373800 582200 374400
rect 576800 371800 582200 372400
rect 576800 369800 582200 370400
rect 475800 256000 477200 257400
rect 475800 254000 477200 255400
rect 475800 252000 477200 253400
rect 475800 250000 477200 251400
rect 475800 248000 477200 249400
rect 475800 246000 477200 247400
rect 475800 244000 477200 245400
rect 475800 242000 477200 243400
rect 475800 240000 477200 241400
rect 568700 241520 569770 241530
rect 568700 240400 577420 241520
rect 568700 240370 576370 240400
rect 475800 238000 477200 239400
rect 475800 236000 477200 237400
rect 475800 234000 477200 235400
rect 475800 232000 477200 233400
rect 475800 230000 477200 231400
rect 475800 228000 477200 229400
rect 475800 226000 477200 227400
rect 475800 224000 477200 225400
rect 475800 222000 477200 223400
rect 475800 220000 477200 221400
rect 475800 218000 477200 219400
rect 475800 216000 477200 217400
rect 475800 214000 477200 215400
rect 475800 212000 477200 213400
rect 475800 210000 477200 211400
rect 475800 208000 477200 209400
rect 475800 206000 477200 207400
rect 475800 204000 477200 205400
rect 475800 202000 477200 203400
rect 475800 200000 477200 201400
rect 475800 198000 477200 199400
rect 475800 196000 477200 197400
rect 475800 194000 477200 195400
rect 475800 192000 477200 193400
rect 475800 190000 477200 191400
rect 579460 198160 580960 201000
rect 579500 189900 580900 198160
rect 475800 188000 477200 189400
rect 475800 186000 477200 187400
rect 475800 184000 477200 185400
rect 475800 182000 477200 183400
rect 475800 180000 477200 181400
rect 475800 178000 477200 179400
rect 475800 176000 477200 177400
rect 475800 174000 477200 175400
rect 475800 172000 477200 173400
rect 475800 170000 477200 171400
rect 475800 168000 477200 169400
rect 475800 166000 477200 167400
rect 576400 167200 579400 175500
rect 475800 164000 477200 165400
rect 475800 162000 477200 163400
rect 475800 160000 477200 161400
rect 475800 158000 477200 159400
rect 475800 156000 477200 157400
rect 475800 154000 477200 155400
rect 475800 152000 477200 153400
rect 475800 150000 477200 151400
rect 475800 148000 477200 149400
rect 475800 146000 477200 147400
rect 475800 144000 477200 145400
rect 475800 142000 477200 143400
rect 573200 151830 576200 152000
rect 573150 148990 576200 151830
rect 573200 143700 576200 148990
rect 475800 140000 477200 141400
rect 475800 138000 477200 139400
rect 475800 136000 477200 137400
rect 475800 134000 477200 135400
rect 475800 132000 477200 133400
rect 475800 130000 477200 131400
rect 475800 128000 477200 129400
rect 475800 126000 477200 127400
rect 475800 124000 477200 125400
rect 475800 122000 477200 123400
rect 570850 123430 570900 130770
rect 570900 123430 577320 130770
rect 570850 123400 577320 123430
rect 475800 120000 477200 121400
rect 475800 118000 477200 119400
rect 475800 116000 477200 117400
rect 475800 114000 477200 115400
rect 475800 112000 477200 113400
rect 475800 110000 477200 111400
rect 475800 108000 477200 109400
rect 475800 106000 477200 107400
rect 475800 104000 477200 105400
rect 475800 102000 477200 103400
rect 475800 100000 477200 101400
rect 475800 98000 477200 99400
rect 475800 96000 477200 97400
rect 475800 94000 477200 95400
rect 475800 92000 477200 93400
rect 475800 90000 477200 91400
rect 475800 88000 477200 89400
rect 475800 86000 477200 87400
rect 475800 84000 477200 85400
rect 475800 82000 477200 83400
rect 475800 80000 477200 81400
rect 475800 78000 477200 79400
rect 475800 76000 477200 77400
rect 475800 74000 477200 75400
rect 475800 72000 477200 73400
rect 475800 70000 477200 71400
rect 475800 68000 477200 69400
rect 475800 66000 477200 67400
rect 475800 64000 477200 65400
rect 475800 62000 477200 63400
rect 475800 60000 477200 61400
rect 475800 58000 477200 59400
rect 475800 56000 477200 57400
rect 475800 54000 477200 55400
rect 475800 52000 477200 53400
rect 475800 50000 477200 51400
rect 475800 48000 477200 49400
rect 475800 46000 477200 47400
rect 475800 44000 477200 45400
rect 475800 42000 477200 43400
rect 475800 40000 477200 41400
rect 475800 38000 477200 39400
rect 475800 36000 477200 37400
rect 475800 34000 477200 35400
rect 475800 32000 477200 33400
rect 475800 30000 477200 31400
rect 475800 28000 477200 29400
rect 475800 26000 477200 27400
rect 475800 24000 477200 25400
rect 475800 22000 477200 23400
rect 475800 20000 477200 21400
rect 475800 18000 477200 19400
rect 475800 16000 477200 17400
rect 475800 14000 477200 15400
rect 475800 12000 477200 13400
rect 475800 10000 477200 11400
rect 475800 8000 477200 9400
rect 475800 6000 477200 7400
rect 475800 4000 477200 5400
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702990 232594 704800
rect 227594 702520 233090 702990
rect 227594 702300 228670 702520
rect 228240 701850 228670 702300
rect 232530 701850 233090 702520
rect 318994 702300 323994 704800
rect 329294 702880 334294 704800
rect 510600 703440 525450 703780
rect 329294 702410 334900 702880
rect 329294 702300 330480 702410
rect 228240 701380 233090 701850
rect 330050 701740 330480 702300
rect 334340 701740 334900 702410
rect 330050 701270 334900 701740
rect 222200 698800 227200 699600
rect 222200 698000 222600 698800
rect 226600 698000 227200 698800
rect 222200 697600 227200 698000
rect 222200 696800 222600 697600
rect 226600 696800 227200 697600
rect 222200 696400 227200 696800
rect 222200 695600 222600 696400
rect 226600 695600 227200 696400
rect 222200 694400 227200 695600
rect 323800 698800 328800 699600
rect 323800 698000 324200 698800
rect 328200 698000 328800 698800
rect 323800 697600 328800 698000
rect 323800 696800 324200 697600
rect 328200 696800 328800 697600
rect 323800 696400 328800 696800
rect 323800 695600 324200 696400
rect 328200 695600 328800 696400
rect 510600 696600 510880 703440
rect 525130 696600 525450 703440
rect 510600 696230 525450 696600
rect 323800 694400 328800 695600
rect 550800 694400 566600 694600
rect 3800 691800 566600 694400
rect 3800 691600 535600 691800
rect 3800 690200 7200 691600
rect 9000 690200 11000 691600
rect 12800 691400 535600 691600
rect 12800 690200 15800 691400
rect 16800 690200 18800 691400
rect 19800 690200 21800 691400
rect 22800 690200 24800 691400
rect 25800 690200 27800 691400
rect 28800 690200 30800 691400
rect 31800 690200 33800 691400
rect 34800 690200 36800 691400
rect 37800 690200 39800 691400
rect 40800 690200 42800 691400
rect 43800 690200 45800 691400
rect 46800 690200 48800 691400
rect 49800 690200 51800 691400
rect 52800 690200 54800 691400
rect 55800 690200 57800 691400
rect 58800 690200 60800 691400
rect 61800 690200 63800 691400
rect 64800 690200 66800 691400
rect 67800 690200 69800 691400
rect 70800 690200 72800 691400
rect 73800 690200 75800 691400
rect 76800 690200 78800 691400
rect 79800 690200 81800 691400
rect 82800 690200 84800 691400
rect 85800 690200 87800 691400
rect 88800 690200 90800 691400
rect 91800 690200 93800 691400
rect 94800 690200 96800 691400
rect 97800 690200 99800 691400
rect 100800 690200 102800 691400
rect 103800 690200 105800 691400
rect 106800 690200 108800 691400
rect 109800 690200 111800 691400
rect 112800 690200 114800 691400
rect 115800 690200 117800 691400
rect 118800 690200 120800 691400
rect 121800 690200 123800 691400
rect 124800 690200 126800 691400
rect 127800 690200 129800 691400
rect 130800 690200 132800 691400
rect 133800 690200 135800 691400
rect 136800 690200 138800 691400
rect 139800 690200 141800 691400
rect 142800 690200 144800 691400
rect 145800 690200 147800 691400
rect 148800 690200 150800 691400
rect 151800 690200 153800 691400
rect 154800 690200 156800 691400
rect 157800 690200 159800 691400
rect 160800 690200 162800 691400
rect 163800 690200 165800 691400
rect 166800 690200 168800 691400
rect 169800 690200 171800 691400
rect 172800 690200 174800 691400
rect 175800 690200 177800 691400
rect 178800 690200 180800 691400
rect 181800 690200 183800 691400
rect 184800 690200 186800 691400
rect 187800 690200 189800 691400
rect 190800 690200 192800 691400
rect 193800 690200 195800 691400
rect 196800 690200 198800 691400
rect 199800 690200 201800 691400
rect 202800 690200 204800 691400
rect 205800 690200 207800 691400
rect 208800 690200 210800 691400
rect 211800 690200 213800 691400
rect 214800 690200 216800 691400
rect 217800 690200 219800 691400
rect 220800 690200 222800 691400
rect 223800 690200 225800 691400
rect 226800 690200 228800 691400
rect 229800 690200 231800 691400
rect 232800 690200 234800 691400
rect 235800 690200 237800 691400
rect 238800 690200 240800 691400
rect 241800 690200 243800 691400
rect 244800 690200 246800 691400
rect 247800 690200 249800 691400
rect 250800 690200 252800 691400
rect 253800 690200 255800 691400
rect 256800 690200 258800 691400
rect 259800 690200 261800 691400
rect 262800 690200 264800 691400
rect 265800 690200 267800 691400
rect 268800 690200 270800 691400
rect 271800 690200 273800 691400
rect 274800 690200 276800 691400
rect 277800 690200 279800 691400
rect 280800 690200 282800 691400
rect 283800 690200 285800 691400
rect 286800 690200 288800 691400
rect 289800 690200 291800 691400
rect 292800 690200 294800 691400
rect 295800 690200 297800 691400
rect 298800 690200 300800 691400
rect 301800 690200 303800 691400
rect 304800 690200 306800 691400
rect 307800 690200 309800 691400
rect 310800 690200 312800 691400
rect 313800 690200 315800 691400
rect 316800 690200 318800 691400
rect 319800 690200 321800 691400
rect 322800 690200 324800 691400
rect 325800 690200 327800 691400
rect 328800 690200 330800 691400
rect 331800 690200 333800 691400
rect 334800 690200 336800 691400
rect 337800 690200 339800 691400
rect 340800 690200 342800 691400
rect 343800 690200 345800 691400
rect 346800 690200 348800 691400
rect 349800 690200 351800 691400
rect 352800 690200 354800 691400
rect 355800 690200 357800 691400
rect 358800 690200 360800 691400
rect 361800 690200 363800 691400
rect 364800 690200 366800 691400
rect 367800 690200 369800 691400
rect 370800 690200 372800 691400
rect 373800 690200 375800 691400
rect 376800 690200 378800 691400
rect 379800 690200 381800 691400
rect 382800 690200 384800 691400
rect 385800 690200 387800 691400
rect 388800 690200 390800 691400
rect 391800 690200 393800 691400
rect 394800 690200 396800 691400
rect 397800 690200 399800 691400
rect 400800 690200 402800 691400
rect 403800 690200 405800 691400
rect 406800 690200 408800 691400
rect 409800 690200 411800 691400
rect 412800 690200 414800 691400
rect 415800 690200 417800 691400
rect 418800 690200 420800 691400
rect 421800 690200 423800 691400
rect 424800 690200 426800 691400
rect 427800 690200 429800 691400
rect 430800 690200 432800 691400
rect 433800 690200 435800 691400
rect 436800 690200 438800 691400
rect 439800 690200 441800 691400
rect 442800 690200 444800 691400
rect 445800 690200 447800 691400
rect 448800 690200 450800 691400
rect 451800 690200 453800 691400
rect 454800 690200 456800 691400
rect 457800 690200 459800 691400
rect 460800 690200 462800 691400
rect 463800 690200 465800 691400
rect 466800 690200 468800 691400
rect 469800 690200 471800 691400
rect 472800 690200 474800 691400
rect 475800 690200 477800 691400
rect 478800 690200 480800 691400
rect 481800 690200 483800 691400
rect 484800 690200 486800 691400
rect 487800 690200 489800 691400
rect 490800 690200 492800 691400
rect 493800 690200 495800 691400
rect 496800 690200 498800 691400
rect 499800 690200 501800 691400
rect 502800 690200 504800 691400
rect 505800 690200 507800 691400
rect 508800 690200 510800 691400
rect 511800 690200 513800 691400
rect 514800 690200 516800 691400
rect 517800 690200 519800 691400
rect 520800 690200 522800 691400
rect 523800 690200 525800 691400
rect 526800 690200 528800 691400
rect 529800 690200 531800 691400
rect 532800 690200 535600 691400
rect 3800 689800 535600 690200
rect 544200 689800 545600 691800
rect 554200 689800 566600 691800
rect 3800 688600 566600 689800
rect 3800 687200 7200 688600
rect 9000 687200 11000 688600
rect 12800 688400 566600 688600
rect 12800 687200 15800 688400
rect 16800 687200 18800 688400
rect 19800 687200 21800 688400
rect 22800 687200 24800 688400
rect 25800 687200 27800 688400
rect 28800 687200 30800 688400
rect 31800 687200 33800 688400
rect 34800 687200 36800 688400
rect 37800 687200 39800 688400
rect 40800 687200 42800 688400
rect 43800 687200 45800 688400
rect 46800 687200 48800 688400
rect 49800 687200 51800 688400
rect 52800 687200 54800 688400
rect 55800 687200 57800 688400
rect 58800 687200 60800 688400
rect 61800 687200 63800 688400
rect 64800 687200 66800 688400
rect 67800 687200 69800 688400
rect 70800 687200 72800 688400
rect 73800 687200 75800 688400
rect 76800 687200 78800 688400
rect 79800 687200 81800 688400
rect 82800 687200 84800 688400
rect 85800 687200 87800 688400
rect 88800 687200 90800 688400
rect 91800 687200 93800 688400
rect 94800 687200 96800 688400
rect 97800 687200 99800 688400
rect 100800 687200 102800 688400
rect 103800 687200 105800 688400
rect 106800 687200 108800 688400
rect 109800 687200 111800 688400
rect 112800 687200 114800 688400
rect 115800 687200 117800 688400
rect 118800 687200 120800 688400
rect 121800 687200 123800 688400
rect 124800 687200 126800 688400
rect 127800 687200 129800 688400
rect 130800 687200 132800 688400
rect 133800 687200 135800 688400
rect 136800 687200 138800 688400
rect 139800 687200 141800 688400
rect 142800 687200 144800 688400
rect 145800 687200 147800 688400
rect 148800 687200 150800 688400
rect 151800 687200 153800 688400
rect 154800 687200 156800 688400
rect 157800 687200 159800 688400
rect 160800 687200 162800 688400
rect 163800 687200 165800 688400
rect 166800 687200 168800 688400
rect 169800 687200 171800 688400
rect 172800 687200 174800 688400
rect 175800 687200 177800 688400
rect 178800 687200 180800 688400
rect 181800 687200 183800 688400
rect 184800 687200 186800 688400
rect 187800 687200 189800 688400
rect 190800 687200 192800 688400
rect 193800 687200 195800 688400
rect 196800 687200 198800 688400
rect 199800 687200 201800 688400
rect 202800 687200 204800 688400
rect 205800 687200 207800 688400
rect 208800 687200 210800 688400
rect 211800 687200 213800 688400
rect 214800 687200 216800 688400
rect 217800 687200 219800 688400
rect 220800 687200 222800 688400
rect 223800 687200 225800 688400
rect 226800 687200 228800 688400
rect 229800 687200 231800 688400
rect 232800 687200 234800 688400
rect 235800 687200 237800 688400
rect 238800 687200 240800 688400
rect 241800 687200 243800 688400
rect 244800 687200 246800 688400
rect 247800 687200 249800 688400
rect 250800 687200 252800 688400
rect 253800 687200 255800 688400
rect 256800 687200 258800 688400
rect 259800 687200 261800 688400
rect 262800 687200 264800 688400
rect 265800 687200 267800 688400
rect 268800 687200 270800 688400
rect 271800 687200 273800 688400
rect 274800 687200 276800 688400
rect 277800 687200 279800 688400
rect 280800 687200 282800 688400
rect 283800 687200 285800 688400
rect 286800 687200 288800 688400
rect 289800 687200 291800 688400
rect 292800 687200 294800 688400
rect 295800 687200 297800 688400
rect 298800 687200 300800 688400
rect 301800 687200 303800 688400
rect 304800 687200 306800 688400
rect 307800 687200 309800 688400
rect 310800 687200 312800 688400
rect 313800 687200 315800 688400
rect 316800 687200 318800 688400
rect 319800 687200 321800 688400
rect 322800 687200 324800 688400
rect 325800 687200 327800 688400
rect 328800 687200 330800 688400
rect 331800 687200 333800 688400
rect 334800 687200 336800 688400
rect 337800 687200 339800 688400
rect 340800 687200 342800 688400
rect 343800 687200 345800 688400
rect 346800 687200 348800 688400
rect 349800 687200 351800 688400
rect 352800 687200 354800 688400
rect 355800 687200 357800 688400
rect 358800 687200 360800 688400
rect 361800 687200 363800 688400
rect 364800 687200 366800 688400
rect 367800 687200 369800 688400
rect 370800 687200 372800 688400
rect 373800 687200 375800 688400
rect 376800 687200 378800 688400
rect 379800 687200 381800 688400
rect 382800 687200 384800 688400
rect 385800 687200 387800 688400
rect 388800 687200 390800 688400
rect 391800 687200 393800 688400
rect 394800 687200 396800 688400
rect 397800 687200 399800 688400
rect 400800 687200 402800 688400
rect 403800 687200 405800 688400
rect 406800 687200 408800 688400
rect 409800 687200 411800 688400
rect 412800 687200 414800 688400
rect 415800 687200 417800 688400
rect 418800 687200 420800 688400
rect 421800 687200 423800 688400
rect 424800 687200 426800 688400
rect 427800 687200 429800 688400
rect 430800 687200 432800 688400
rect 433800 687200 435800 688400
rect 436800 687200 438800 688400
rect 439800 687200 441800 688400
rect 442800 687200 444800 688400
rect 445800 687200 447800 688400
rect 448800 687200 450800 688400
rect 451800 687200 453800 688400
rect 454800 687200 456800 688400
rect 457800 687200 459800 688400
rect 460800 687200 462800 688400
rect 463800 687200 465800 688400
rect 466800 687200 468800 688400
rect 469800 687200 471800 688400
rect 472800 687200 474800 688400
rect 475800 687200 477800 688400
rect 478800 687200 480800 688400
rect 481800 687200 483800 688400
rect 484800 687200 486800 688400
rect 487800 687200 489800 688400
rect 490800 687200 492800 688400
rect 493800 687200 495800 688400
rect 496800 687200 498800 688400
rect 499800 687200 501800 688400
rect 502800 687200 504800 688400
rect 505800 687200 507800 688400
rect 508800 687200 510800 688400
rect 511800 687200 513800 688400
rect 514800 687200 516800 688400
rect 517800 687200 519800 688400
rect 520800 687200 522800 688400
rect 523800 687200 525800 688400
rect 526800 687200 528800 688400
rect 529800 687200 531800 688400
rect 532800 687800 566600 688400
rect 532800 687200 535600 687800
rect 3800 685800 535600 687200
rect 544200 685800 545600 687800
rect 554200 685800 566600 687800
rect 3800 685600 566600 685800
rect 3800 684200 7200 685600
rect 9000 684200 11000 685600
rect 12800 685400 566600 685600
rect 12800 684200 15800 685400
rect 16800 684200 18800 685400
rect 19800 684200 21800 685400
rect 22800 684200 24800 685400
rect 25800 684200 27800 685400
rect 28800 684200 30800 685400
rect 31800 684200 33800 685400
rect 34800 684200 36800 685400
rect 37800 684200 39800 685400
rect 40800 684200 42800 685400
rect 43800 684200 45800 685400
rect 46800 684200 48800 685400
rect 49800 684200 51800 685400
rect 52800 684200 54800 685400
rect 55800 684200 57800 685400
rect 58800 684200 60800 685400
rect 61800 684200 63800 685400
rect 64800 684200 66800 685400
rect 67800 684200 69800 685400
rect 70800 684200 72800 685400
rect 73800 684200 75800 685400
rect 76800 684200 78800 685400
rect 79800 684200 81800 685400
rect 82800 684200 84800 685400
rect 85800 684200 87800 685400
rect 88800 684200 90800 685400
rect 91800 684200 93800 685400
rect 94800 684200 96800 685400
rect 97800 684200 99800 685400
rect 100800 684200 102800 685400
rect 103800 684200 105800 685400
rect 106800 684200 108800 685400
rect 109800 684200 111800 685400
rect 112800 684200 114800 685400
rect 115800 684200 117800 685400
rect 118800 684200 120800 685400
rect 121800 684200 123800 685400
rect 124800 684200 126800 685400
rect 127800 684200 129800 685400
rect 130800 684200 132800 685400
rect 133800 684200 135800 685400
rect 136800 684200 138800 685400
rect 139800 684200 141800 685400
rect 142800 684200 144800 685400
rect 145800 684200 147800 685400
rect 148800 684200 150800 685400
rect 151800 684200 153800 685400
rect 154800 684200 156800 685400
rect 157800 684200 159800 685400
rect 160800 684200 162800 685400
rect 163800 684200 165800 685400
rect 166800 684200 168800 685400
rect 169800 684200 171800 685400
rect 172800 684200 174800 685400
rect 175800 684200 177800 685400
rect 178800 684200 180800 685400
rect 181800 684200 183800 685400
rect 184800 684200 186800 685400
rect 187800 684200 189800 685400
rect 190800 684200 192800 685400
rect 193800 684200 195800 685400
rect 196800 684200 198800 685400
rect 199800 684200 201800 685400
rect 202800 684200 204800 685400
rect 205800 684200 207800 685400
rect 208800 684200 210800 685400
rect 211800 684200 213800 685400
rect 214800 684200 216800 685400
rect 217800 684200 219800 685400
rect 220800 684200 222800 685400
rect 223800 684200 225800 685400
rect 226800 684200 228800 685400
rect 229800 684200 231800 685400
rect 232800 684200 234800 685400
rect 235800 684200 237800 685400
rect 238800 684200 240800 685400
rect 241800 684200 243800 685400
rect 244800 684200 246800 685400
rect 247800 684200 249800 685400
rect 250800 684200 252800 685400
rect 253800 684200 255800 685400
rect 256800 684200 258800 685400
rect 259800 684200 261800 685400
rect 262800 684200 264800 685400
rect 265800 684200 267800 685400
rect 268800 684200 270800 685400
rect 271800 684200 273800 685400
rect 274800 684200 276800 685400
rect 277800 684200 279800 685400
rect 280800 684200 282800 685400
rect 283800 684200 285800 685400
rect 286800 684200 288800 685400
rect 289800 684200 291800 685400
rect 292800 684200 294800 685400
rect 295800 684200 297800 685400
rect 298800 684200 300800 685400
rect 301800 684200 303800 685400
rect 304800 684200 306800 685400
rect 307800 684200 309800 685400
rect 310800 684200 312800 685400
rect 313800 684200 315800 685400
rect 316800 684200 318800 685400
rect 319800 684200 321800 685400
rect 322800 684200 324800 685400
rect 325800 684200 327800 685400
rect 328800 684200 330800 685400
rect 331800 684200 333800 685400
rect 334800 684200 336800 685400
rect 337800 684200 339800 685400
rect 340800 684200 342800 685400
rect 343800 684200 345800 685400
rect 346800 684200 348800 685400
rect 349800 684200 351800 685400
rect 352800 684200 354800 685400
rect 355800 684200 357800 685400
rect 358800 684200 360800 685400
rect 361800 684200 363800 685400
rect 364800 684200 366800 685400
rect 367800 684200 369800 685400
rect 370800 684200 372800 685400
rect 373800 684200 375800 685400
rect 376800 684200 378800 685400
rect 379800 684200 381800 685400
rect 382800 684200 384800 685400
rect 385800 684200 387800 685400
rect 388800 684200 390800 685400
rect 391800 684200 393800 685400
rect 394800 684200 396800 685400
rect 397800 684200 399800 685400
rect 400800 684200 402800 685400
rect 403800 684200 405800 685400
rect 406800 684200 408800 685400
rect 409800 684200 411800 685400
rect 412800 684200 414800 685400
rect 415800 684200 417800 685400
rect 418800 684200 420800 685400
rect 421800 684200 423800 685400
rect 424800 684200 426800 685400
rect 427800 684200 429800 685400
rect 430800 684200 432800 685400
rect 433800 684200 435800 685400
rect 436800 684200 438800 685400
rect 439800 684200 441800 685400
rect 442800 684200 444800 685400
rect 445800 684200 447800 685400
rect 448800 684200 450800 685400
rect 451800 684200 453800 685400
rect 454800 684200 456800 685400
rect 457800 684200 459800 685400
rect 460800 684200 462800 685400
rect 463800 684200 465800 685400
rect 466800 684200 468800 685400
rect 469800 684200 471800 685400
rect 472800 684200 474800 685400
rect 475800 684200 477800 685400
rect 478800 684200 480800 685400
rect 481800 684200 483800 685400
rect 484800 684200 486800 685400
rect 487800 684200 489800 685400
rect 490800 684200 492800 685400
rect 493800 684200 495800 685400
rect 496800 684200 498800 685400
rect 499800 684200 501800 685400
rect 502800 684200 504800 685400
rect 505800 684200 507800 685400
rect 508800 684200 510800 685400
rect 511800 684200 513800 685400
rect 514800 684200 516800 685400
rect 517800 684200 519800 685400
rect 520800 684200 522800 685400
rect 523800 684200 525800 685400
rect 526800 684200 528800 685400
rect 529800 684200 531800 685400
rect 532800 684200 566600 685400
rect 3800 683800 566600 684200
rect 3800 682600 535600 683800
rect 3800 681200 7200 682600
rect 9000 681200 11000 682600
rect 12800 682400 535600 682600
rect 12800 681200 15800 682400
rect 16800 681200 18800 682400
rect 19800 681200 21800 682400
rect 22800 681200 24800 682400
rect 25800 681200 27800 682400
rect 28800 681200 30800 682400
rect 31800 681200 33800 682400
rect 34800 681200 36800 682400
rect 37800 681200 39800 682400
rect 40800 681200 42800 682400
rect 43800 681200 45800 682400
rect 46800 681200 48800 682400
rect 49800 681200 51800 682400
rect 52800 681200 54800 682400
rect 55800 681200 57800 682400
rect 58800 681200 60800 682400
rect 61800 681200 63800 682400
rect 64800 681200 66800 682400
rect 67800 681200 69800 682400
rect 70800 681200 72800 682400
rect 73800 681200 75800 682400
rect 76800 681200 78800 682400
rect 79800 681200 81800 682400
rect 82800 681200 84800 682400
rect 85800 681200 87800 682400
rect 88800 681200 90800 682400
rect 91800 681200 93800 682400
rect 94800 681200 96800 682400
rect 97800 681200 99800 682400
rect 100800 681200 102800 682400
rect 103800 681200 105800 682400
rect 106800 681200 108800 682400
rect 109800 681200 111800 682400
rect 112800 681200 114800 682400
rect 115800 681200 117800 682400
rect 118800 681200 120800 682400
rect 121800 681200 123800 682400
rect 124800 681200 126800 682400
rect 127800 681200 129800 682400
rect 130800 681200 132800 682400
rect 133800 681200 135800 682400
rect 136800 681200 138800 682400
rect 139800 681200 141800 682400
rect 142800 681200 144800 682400
rect 145800 681200 147800 682400
rect 148800 681200 150800 682400
rect 151800 681200 153800 682400
rect 154800 681200 156800 682400
rect 157800 681200 159800 682400
rect 160800 681200 162800 682400
rect 163800 681200 165800 682400
rect 166800 681200 168800 682400
rect 169800 681200 171800 682400
rect 172800 681200 174800 682400
rect 175800 681200 177800 682400
rect 178800 681200 180800 682400
rect 181800 681200 183800 682400
rect 184800 681200 186800 682400
rect 187800 681200 189800 682400
rect 190800 681200 192800 682400
rect 193800 681200 195800 682400
rect 196800 681200 198800 682400
rect 199800 681200 201800 682400
rect 202800 681200 204800 682400
rect 205800 681200 207800 682400
rect 208800 681200 210800 682400
rect 211800 681200 213800 682400
rect 214800 681200 216800 682400
rect 217800 681200 219800 682400
rect 220800 681200 222800 682400
rect 223800 681200 225800 682400
rect 226800 681200 228800 682400
rect 229800 681200 231800 682400
rect 232800 681200 234800 682400
rect 235800 681200 237800 682400
rect 238800 681200 240800 682400
rect 241800 681200 243800 682400
rect 244800 681200 246800 682400
rect 247800 681200 249800 682400
rect 250800 681200 252800 682400
rect 253800 681200 255800 682400
rect 256800 681200 258800 682400
rect 259800 681200 261800 682400
rect 262800 681200 264800 682400
rect 265800 681200 267800 682400
rect 268800 681200 270800 682400
rect 271800 681200 273800 682400
rect 274800 681200 276800 682400
rect 277800 681200 279800 682400
rect 280800 681200 282800 682400
rect 283800 681200 285800 682400
rect 286800 681200 288800 682400
rect 289800 681200 291800 682400
rect 292800 681200 294800 682400
rect 295800 681200 297800 682400
rect 298800 681200 300800 682400
rect 301800 681200 303800 682400
rect 304800 681200 306800 682400
rect 307800 681200 309800 682400
rect 310800 681200 312800 682400
rect 313800 681200 315800 682400
rect 316800 681200 318800 682400
rect 319800 681200 321800 682400
rect 322800 681200 324800 682400
rect 325800 681200 327800 682400
rect 328800 681200 330800 682400
rect 331800 681200 333800 682400
rect 334800 681200 336800 682400
rect 337800 681200 339800 682400
rect 340800 681200 342800 682400
rect 343800 681200 345800 682400
rect 346800 681200 348800 682400
rect 349800 681200 351800 682400
rect 352800 681200 354800 682400
rect 355800 681200 357800 682400
rect 358800 681200 360800 682400
rect 361800 681200 363800 682400
rect 364800 681200 366800 682400
rect 367800 681200 369800 682400
rect 370800 681200 372800 682400
rect 373800 681200 375800 682400
rect 376800 681200 378800 682400
rect 379800 681200 381800 682400
rect 382800 681200 384800 682400
rect 385800 681200 387800 682400
rect 388800 681200 390800 682400
rect 391800 681200 393800 682400
rect 394800 681200 396800 682400
rect 397800 681200 399800 682400
rect 400800 681200 402800 682400
rect 403800 681200 405800 682400
rect 406800 681200 408800 682400
rect 409800 681200 411800 682400
rect 412800 681200 414800 682400
rect 415800 681200 417800 682400
rect 418800 681200 420800 682400
rect 421800 681200 423800 682400
rect 424800 681200 426800 682400
rect 427800 681200 429800 682400
rect 430800 681200 432800 682400
rect 433800 681200 435800 682400
rect 436800 681200 438800 682400
rect 439800 681200 441800 682400
rect 442800 681200 444800 682400
rect 445800 681200 447800 682400
rect 448800 681200 450800 682400
rect 451800 681200 453800 682400
rect 454800 681200 456800 682400
rect 457800 681200 459800 682400
rect 460800 681200 462800 682400
rect 463800 681200 465800 682400
rect 466800 681200 468800 682400
rect 469800 681200 471800 682400
rect 472800 681200 474800 682400
rect 475800 681200 477800 682400
rect 478800 681200 480800 682400
rect 481800 681200 483800 682400
rect 484800 681200 486800 682400
rect 487800 681200 489800 682400
rect 490800 681200 492800 682400
rect 493800 681200 495800 682400
rect 496800 681200 498800 682400
rect 499800 681200 501800 682400
rect 502800 681200 504800 682400
rect 505800 681200 507800 682400
rect 508800 681200 510800 682400
rect 511800 681200 513800 682400
rect 514800 681200 516800 682400
rect 517800 681200 519800 682400
rect 520800 681200 522800 682400
rect 523800 681200 525800 682400
rect 526800 681200 528800 682400
rect 529800 681200 531800 682400
rect 532800 681800 535600 682400
rect 544200 681800 545600 683800
rect 554200 681800 566600 683800
rect 532800 681200 566600 681800
rect 3800 679800 566600 681200
rect 3800 679600 535600 679800
rect 3800 678200 7200 679600
rect 9000 678200 11000 679600
rect 12800 678200 15000 679600
rect 3800 676600 15000 678200
rect 3800 675200 7200 676600
rect 9000 675200 11000 676600
rect 12800 675200 15000 676600
rect 3800 673600 15000 675200
rect 3800 672200 7200 673600
rect 9000 672200 11000 673600
rect 12800 672200 15000 673600
rect 3800 670600 15000 672200
rect 3800 669200 7200 670600
rect 9000 669200 11000 670600
rect 12800 669200 15000 670600
rect 3800 667600 15000 669200
rect 3800 666200 7200 667600
rect 9000 666200 11000 667600
rect 12800 666200 15000 667600
rect 3800 664600 15000 666200
rect 3800 663200 7200 664600
rect 9000 663200 11000 664600
rect 12800 663200 15000 664600
rect 3800 661600 15000 663200
rect 3800 660200 7200 661600
rect 9000 660200 11000 661600
rect 12800 660200 15000 661600
rect 3800 658600 15000 660200
rect 3800 657200 7200 658600
rect 9000 657200 11000 658600
rect 12800 657200 15000 658600
rect 3800 656000 15000 657200
rect 3800 654800 4800 656000
rect 6200 655600 15000 656000
rect 6200 654800 7200 655600
rect 3800 654200 7200 654800
rect 9000 654200 11000 655600
rect 12800 654200 15000 655600
rect 3800 654000 15000 654200
rect 3800 653800 4800 654000
rect 600 652800 4800 653800
rect 6200 652800 15000 654000
rect 600 652600 15000 652800
rect 600 652000 7200 652600
rect 600 650800 4800 652000
rect 6200 651200 7200 652000
rect 9000 651200 11000 652600
rect 12800 651200 15000 652600
rect 6200 650800 15000 651200
rect 600 650000 15000 650800
rect 600 649600 4800 650000
rect 200 648800 4800 649600
rect 6200 649600 15000 650000
rect 6200 648800 7200 649600
rect 200 648200 7200 648800
rect 9000 648200 11000 649600
rect 12800 648200 15000 649600
rect 200 648000 15000 648200
rect 200 646800 4800 648000
rect 6200 646800 15000 648000
rect 200 646600 15000 646800
rect 200 646000 7200 646600
rect 200 644800 4800 646000
rect 6200 645200 7200 646000
rect 9000 645200 11000 646600
rect 12800 645200 15000 646600
rect 6200 644800 15000 645200
rect 200 644000 15000 644800
rect 200 642800 4800 644000
rect 6200 643600 15000 644000
rect 6200 642800 7200 643600
rect 200 642200 7200 642800
rect 9000 642200 11000 643600
rect 12800 642200 15000 643600
rect 200 642000 15000 642200
rect 200 640800 4800 642000
rect 6200 640800 15000 642000
rect 200 640600 15000 640800
rect 200 640000 7200 640600
rect 200 638800 4800 640000
rect 6200 639200 7200 640000
rect 9000 639200 11000 640600
rect 12800 639200 15000 640600
rect 6200 638800 15000 639200
rect 200 638000 15000 638800
rect 200 636800 4800 638000
rect 6200 637600 15000 638000
rect 6200 636800 7200 637600
rect 200 636200 7200 636800
rect 9000 636200 11000 637600
rect 12800 636200 15000 637600
rect 200 636000 15000 636200
rect 200 634800 4800 636000
rect 6200 634800 15000 636000
rect 200 634600 15000 634800
rect 200 634000 7200 634600
rect 200 633200 4800 634000
rect 600 632800 4800 633200
rect 6200 633200 7200 634000
rect 9000 633200 11000 634600
rect 12800 633200 15000 634600
rect 6200 632800 15000 633200
rect 600 632000 15000 632800
rect 600 631800 4800 632000
rect 4400 630800 4800 631800
rect 6200 630800 7400 632000
rect 8800 631800 15000 632000
rect 475200 677400 477800 678200
rect 475200 676000 475800 677400
rect 477200 676000 477800 677400
rect 475200 675400 477800 676000
rect 475200 674000 475800 675400
rect 477200 674000 477800 675400
rect 475200 673400 477800 674000
rect 475200 672000 475800 673400
rect 477200 672000 477800 673400
rect 475200 671400 477800 672000
rect 475200 670000 475800 671400
rect 477200 670000 477800 671400
rect 534800 677800 535600 679600
rect 544200 677800 545600 679800
rect 554200 677800 566600 679800
rect 534800 675800 566600 677800
rect 534800 673800 535600 675800
rect 544200 673800 545600 675800
rect 554200 673800 566600 675800
rect 534800 671800 566600 673800
rect 475200 669400 477800 670000
rect 475200 668000 475800 669400
rect 477200 668000 477800 669400
rect 475200 667400 477800 668000
rect 475200 666000 475800 667400
rect 477200 666000 477800 667400
rect 475200 665400 477800 666000
rect 475200 664000 475800 665400
rect 477200 664000 477800 665400
rect 475200 663400 477800 664000
rect 519680 669740 527080 670340
rect 519680 664340 520580 669740
rect 526480 664340 527080 669740
rect 519680 663640 527080 664340
rect 534800 669800 535600 671800
rect 544200 669800 545600 671800
rect 554200 669800 566600 671800
rect 534800 667800 566600 669800
rect 534800 665800 535600 667800
rect 544200 665800 545600 667800
rect 554200 665800 566600 667800
rect 534800 663800 566600 665800
rect 475200 662000 475800 663400
rect 477200 662000 477800 663400
rect 475200 661400 477800 662000
rect 475200 660000 475800 661400
rect 477200 660000 477800 661400
rect 475200 659400 477800 660000
rect 475200 658000 475800 659400
rect 477200 658000 477800 659400
rect 475200 657400 477800 658000
rect 475200 656000 475800 657400
rect 477200 656000 477800 657400
rect 475200 655400 477800 656000
rect 475200 654000 475800 655400
rect 477200 654000 477800 655400
rect 475200 653400 477800 654000
rect 475200 652000 475800 653400
rect 477200 652000 477800 653400
rect 475200 651400 477800 652000
rect 475200 650000 475800 651400
rect 477200 650000 477800 651400
rect 475200 649400 477800 650000
rect 475200 648000 475800 649400
rect 477200 648000 477800 649400
rect 475200 647400 477800 648000
rect 534800 661800 535600 663800
rect 544200 661800 545600 663800
rect 554200 661800 566600 663800
rect 534800 659800 566600 661800
rect 534800 657800 535600 659800
rect 544200 657800 545600 659800
rect 554200 657800 566600 659800
rect 534800 655800 566600 657800
rect 534800 653800 535600 655800
rect 544200 653800 545600 655800
rect 554200 653800 566600 655800
rect 534800 651800 566600 653800
rect 534800 649800 535600 651800
rect 544200 649800 545600 651800
rect 554200 649800 566600 651800
rect 534800 647800 566600 649800
rect 475200 646000 475800 647400
rect 477200 646000 477800 647400
rect 475200 645400 477800 646000
rect 475200 644000 475800 645400
rect 477200 644000 477800 645400
rect 475200 643400 477800 644000
rect 475200 642000 475800 643400
rect 477200 642000 477800 643400
rect 475200 641400 477800 642000
rect 475200 640000 475800 641400
rect 477200 640000 477800 641400
rect 519780 646740 527180 647440
rect 519780 641340 520780 646740
rect 526680 641340 527180 646740
rect 519780 640740 527180 641340
rect 534800 645800 535600 647800
rect 544200 645800 545600 647800
rect 554200 645800 566600 647800
rect 534800 644400 566600 645800
rect 576350 644400 583900 644590
rect 534800 644270 583900 644400
rect 534800 643800 576690 644270
rect 534800 641800 535600 643800
rect 544200 641800 545600 643800
rect 554200 641800 576690 643800
rect 475200 639400 477800 640000
rect 475200 638000 475800 639400
rect 477200 638000 477800 639400
rect 475200 637400 477800 638000
rect 475200 636000 475800 637400
rect 477200 636000 477800 637400
rect 475200 635400 477800 636000
rect 475200 634000 475800 635400
rect 477200 634000 477800 635400
rect 475200 633400 477800 634000
rect 475200 632000 475800 633400
rect 477200 632000 477800 633400
rect 8800 630800 9200 631800
rect 4400 630000 9200 630800
rect 475200 631400 477800 632000
rect 4400 628800 4800 630000
rect 6200 628800 7400 630000
rect 8800 628800 9200 630000
rect 4400 628000 9200 628800
rect 4400 626800 4800 628000
rect 6200 626800 7400 628000
rect 8800 626800 9200 628000
rect 4400 626000 9200 626800
rect 4400 624800 4800 626000
rect 6200 624800 7400 626000
rect 8800 624800 9200 626000
rect 4400 624000 9200 624800
rect 4400 622800 4800 624000
rect 6200 622800 7400 624000
rect 8800 622800 9200 624000
rect 4400 622000 9200 622800
rect 4400 620800 4800 622000
rect 6200 620800 7400 622000
rect 8800 620800 9200 622000
rect 4400 620000 9200 620800
rect 4400 618800 4800 620000
rect 6200 618800 7400 620000
rect 8800 618800 9200 620000
rect 4400 618000 9200 618800
rect 4400 616800 4800 618000
rect 6200 616800 7400 618000
rect 8800 616800 9200 618000
rect 4400 616000 9200 616800
rect 4400 614800 4800 616000
rect 6200 614800 7400 616000
rect 8800 614800 9200 616000
rect 4400 614000 9200 614800
rect 4400 612800 4800 614000
rect 6200 612800 7400 614000
rect 8800 612800 9200 614000
rect 4400 612000 9200 612800
rect 4400 610800 4800 612000
rect 6200 610800 7400 612000
rect 8800 610800 9200 612000
rect 4400 610000 9200 610800
rect 4400 608800 4800 610000
rect 6200 608800 7400 610000
rect 8800 608800 9200 610000
rect 4400 608000 9200 608800
rect 4400 606800 4800 608000
rect 6200 606800 7400 608000
rect 8800 606800 9200 608000
rect 4400 606000 9200 606800
rect 4400 604800 4800 606000
rect 6200 604800 7400 606000
rect 8800 604800 9200 606000
rect 4400 604000 9200 604800
rect 4400 602800 4800 604000
rect 6200 602800 7400 604000
rect 8800 602800 9200 604000
rect 4400 602000 9200 602800
rect 4400 600800 4800 602000
rect 6200 600800 7400 602000
rect 8800 600800 9200 602000
rect 4400 600000 9200 600800
rect 4400 598800 4800 600000
rect 6200 598800 7400 600000
rect 8800 598800 9200 600000
rect 4400 598000 9200 598800
rect 4400 596800 4800 598000
rect 6200 596800 7400 598000
rect 8800 596800 9200 598000
rect 4400 596000 9200 596800
rect 4400 594800 4800 596000
rect 6200 594800 7400 596000
rect 8800 594800 9200 596000
rect 4400 594000 9200 594800
rect 4400 592800 4800 594000
rect 6200 592800 7400 594000
rect 8800 592800 9200 594000
rect 4400 592000 9200 592800
rect 4400 590800 4800 592000
rect 6200 590800 7400 592000
rect 8800 590800 9200 592000
rect 4400 590000 9200 590800
rect 4400 588800 4800 590000
rect 6200 588800 7400 590000
rect 8800 588800 9200 590000
rect 4400 588000 9200 588800
rect 4400 586800 4800 588000
rect 6200 586800 7400 588000
rect 8800 586800 9200 588000
rect 4400 586000 9200 586800
rect 4400 584800 4800 586000
rect 6200 584800 7400 586000
rect 8800 584800 9200 586000
rect 4400 584000 9200 584800
rect 4400 582800 4800 584000
rect 6200 582800 7400 584000
rect 8800 582800 9200 584000
rect 4400 582000 9200 582800
rect 4400 580800 4800 582000
rect 6200 580800 7400 582000
rect 8800 580800 9200 582000
rect 4400 580000 9200 580800
rect 4400 578800 4800 580000
rect 6200 578800 7400 580000
rect 8800 578800 9200 580000
rect 4400 578000 9200 578800
rect 4400 576800 4800 578000
rect 6200 576800 7400 578000
rect 8800 576800 9200 578000
rect 4400 576000 9200 576800
rect 4400 574800 4800 576000
rect 6200 574800 7400 576000
rect 8800 574800 9200 576000
rect 4400 574000 9200 574800
rect 4400 572800 4800 574000
rect 6200 572800 7400 574000
rect 8800 572800 9200 574000
rect 4400 572000 9200 572800
rect 4400 570800 4800 572000
rect 6200 570800 7400 572000
rect 8800 570800 9200 572000
rect 4400 570000 9200 570800
rect 4400 568800 4800 570000
rect 6200 568800 7400 570000
rect 8800 568800 9200 570000
rect 4400 568000 9200 568800
rect 4400 566800 4800 568000
rect 6200 566800 7400 568000
rect 8800 566800 9200 568000
rect 4400 566000 9200 566800
rect 4400 564800 4800 566000
rect 6200 564800 7400 566000
rect 8800 564800 9200 566000
rect 330 564320 3200 564730
rect 330 549250 870 564320
rect 2600 549250 3200 564320
rect 330 548720 3200 549250
rect 4400 564000 9200 564800
rect 4400 562800 4800 564000
rect 6200 562800 7400 564000
rect 8800 562800 9200 564000
rect 4400 562000 9200 562800
rect 4400 560800 4800 562000
rect 6200 560800 7400 562000
rect 8800 560800 9200 562000
rect 4400 560000 9200 560800
rect 4400 558800 4800 560000
rect 6200 558800 7400 560000
rect 8800 558800 9200 560000
rect 4400 558000 9200 558800
rect 4400 556800 4800 558000
rect 6200 556800 7400 558000
rect 8800 556800 9200 558000
rect 4400 556000 9200 556800
rect 4400 554800 4800 556000
rect 6200 554800 7400 556000
rect 8800 554800 9200 556000
rect 4400 554000 9200 554800
rect 4400 552800 4800 554000
rect 6200 552800 7400 554000
rect 8800 552800 9200 554000
rect 4400 552000 9200 552800
rect 4400 550800 4800 552000
rect 6200 550800 7400 552000
rect 8800 550800 9200 552000
rect 4400 550000 9200 550800
rect 4400 548800 4800 550000
rect 6200 548800 7400 550000
rect 8800 548800 9200 550000
rect 4400 548000 9200 548800
rect 4400 546800 4800 548000
rect 6200 546800 7400 548000
rect 8800 546800 9200 548000
rect 4400 546000 9200 546800
rect 3200 544800 4800 546000
rect 6200 544800 7400 546000
rect 8800 544800 9200 546000
rect 3200 544000 9200 544800
rect 3200 542800 4800 544000
rect 6200 542800 7400 544000
rect 8800 542800 9200 544000
rect 3200 542000 9200 542800
rect 3200 540800 4800 542000
rect 6200 540800 7400 542000
rect 8800 540800 9200 542000
rect 3200 540000 9200 540800
rect 3200 538800 4800 540000
rect 6200 538800 7400 540000
rect 8800 538800 9200 540000
rect 3200 538000 9200 538800
rect 15800 630200 17000 630400
rect 15800 629600 16000 630200
rect 16800 629600 17000 630200
rect 15800 627200 17000 629600
rect 15800 626600 16000 627200
rect 16800 626600 17000 627200
rect 15800 624200 17000 626600
rect 15800 623600 16000 624200
rect 16800 623600 17000 624200
rect 15800 621200 17000 623600
rect 15800 620600 16000 621200
rect 16800 620600 17000 621200
rect 15800 618200 17000 620600
rect 15800 617600 16000 618200
rect 16800 617600 17000 618200
rect 15800 615200 17000 617600
rect 15800 614600 16000 615200
rect 16800 614600 17000 615200
rect 15800 612200 17000 614600
rect 15800 611600 16000 612200
rect 16800 611600 17000 612200
rect 15800 609200 17000 611600
rect 15800 608600 16000 609200
rect 16800 608600 17000 609200
rect 15800 606200 17000 608600
rect 15800 605600 16000 606200
rect 16800 605600 17000 606200
rect 15800 603200 17000 605600
rect 15800 602600 16000 603200
rect 16800 602600 17000 603200
rect 15800 600200 17000 602600
rect 15800 599600 16000 600200
rect 16800 599600 17000 600200
rect 15800 597200 17000 599600
rect 15800 596600 16000 597200
rect 16800 596600 17000 597200
rect 15800 594200 17000 596600
rect 15800 593600 16000 594200
rect 16800 593600 17000 594200
rect 15800 591200 17000 593600
rect 15800 590600 16000 591200
rect 16800 590600 17000 591200
rect 15800 588200 17000 590600
rect 15800 587600 16000 588200
rect 16800 587600 17000 588200
rect 15800 585200 17000 587600
rect 15800 584600 16000 585200
rect 16800 584600 17000 585200
rect 15800 582200 17000 584600
rect 15800 581600 16000 582200
rect 16800 581600 17000 582200
rect 15800 579200 17000 581600
rect 15800 578600 16000 579200
rect 16800 578600 17000 579200
rect 15800 576200 17000 578600
rect 15800 575600 16000 576200
rect 16800 575600 17000 576200
rect 15800 573200 17000 575600
rect 15800 572600 16000 573200
rect 16800 572600 17000 573200
rect 15800 570200 17000 572600
rect 15800 569600 16000 570200
rect 16800 569600 17000 570200
rect 15800 567200 17000 569600
rect 15800 566600 16000 567200
rect 16800 566600 17000 567200
rect 15800 564200 17000 566600
rect 15800 563600 16000 564200
rect 16800 563600 17000 564200
rect 15800 561200 17000 563600
rect 15800 560600 16000 561200
rect 16800 560600 17000 561200
rect 15800 558200 17000 560600
rect 15800 557600 16000 558200
rect 16800 557600 17000 558200
rect 15800 555200 17000 557600
rect 15800 554600 16000 555200
rect 16800 554600 17000 555200
rect 15800 552200 17000 554600
rect 15800 551600 16000 552200
rect 16800 551600 17000 552200
rect 15800 549200 17000 551600
rect 15800 548600 16000 549200
rect 16800 548600 17000 549200
rect 15800 547800 17000 548600
rect 15800 547200 16000 547800
rect 16800 547200 17000 547800
rect 15800 544800 17000 547200
rect 15800 544200 16000 544800
rect 16800 544400 17000 544800
rect 475200 630000 475800 631400
rect 477200 630000 477800 631400
rect 475200 629400 477800 630000
rect 534800 639800 576690 641800
rect 534800 637800 535600 639800
rect 544200 637800 545600 639800
rect 554200 637800 576690 639800
rect 534800 635800 576690 637800
rect 534800 633800 535600 635800
rect 544200 633800 545600 635800
rect 554200 633800 576690 635800
rect 534800 631800 576690 633800
rect 475200 628000 475800 629400
rect 477200 628000 477800 629400
rect 475200 627400 477800 628000
rect 475200 626000 475800 627400
rect 477200 626000 477800 627400
rect 499220 629510 507100 629880
rect 499220 628360 499340 629510
rect 507010 628360 507100 629510
rect 534800 629800 535600 631800
rect 544200 629800 545600 631800
rect 554200 630020 576690 631800
rect 583530 630020 583900 644270
rect 554200 629800 583900 630020
rect 534800 629740 583900 629800
rect 534800 629000 579000 629740
rect 499220 627120 507100 628360
rect 475200 625400 477800 626000
rect 475200 624000 475800 625400
rect 477200 624000 477800 625400
rect 475200 623400 477800 624000
rect 475200 622000 475800 623400
rect 477200 622000 477800 623400
rect 475200 621400 477800 622000
rect 475200 620000 475800 621400
rect 477200 620000 477800 621400
rect 475200 619400 477800 620000
rect 475200 618000 475800 619400
rect 477200 618000 477800 619400
rect 475200 617400 477800 618000
rect 475200 616000 475800 617400
rect 477200 616000 477800 617400
rect 519880 623040 527180 623740
rect 519880 617740 520580 623040
rect 526580 617740 527180 623040
rect 519880 617040 527180 617740
rect 475200 615400 477800 616000
rect 475200 614000 475800 615400
rect 477200 614000 477800 615400
rect 475200 613400 477800 614000
rect 475200 612000 475800 613400
rect 477200 612000 477800 613400
rect 475200 611400 477800 612000
rect 475200 610000 475800 611400
rect 477200 610000 477800 611400
rect 475200 609400 477800 610000
rect 475200 608000 475800 609400
rect 477200 608000 477800 609400
rect 475200 607400 477800 608000
rect 475200 606000 475800 607400
rect 477200 606000 477800 607400
rect 475200 605400 477800 606000
rect 475200 604000 475800 605400
rect 477200 604000 477800 605400
rect 475200 603400 477800 604000
rect 475200 602000 475800 603400
rect 477200 602000 477800 603400
rect 475200 601400 477800 602000
rect 475200 600000 475800 601400
rect 477200 600000 477800 601400
rect 475200 599400 477800 600000
rect 475200 598000 475800 599400
rect 477200 598000 477800 599400
rect 475200 597400 477800 598000
rect 475200 596000 475800 597400
rect 477200 596000 477800 597400
rect 475200 595400 477800 596000
rect 475200 594000 475800 595400
rect 477200 594000 477800 595400
rect 475200 593400 477800 594000
rect 475200 592000 475800 593400
rect 477200 592000 477800 593400
rect 475200 591400 477800 592000
rect 475200 590000 475800 591400
rect 477200 590000 477800 591400
rect 475200 589400 477800 590000
rect 475200 588000 475800 589400
rect 477200 588000 477800 589400
rect 475200 587400 477800 588000
rect 475200 586000 475800 587400
rect 477200 586000 477800 587400
rect 475200 585400 477800 586000
rect 475200 584000 475800 585400
rect 477200 584000 477800 585400
rect 475200 583400 477800 584000
rect 475200 582000 475800 583400
rect 477200 582000 477800 583400
rect 475200 581400 477800 582000
rect 475200 580000 475800 581400
rect 477200 580000 477800 581400
rect 475200 579400 477800 580000
rect 475200 578000 475800 579400
rect 477200 578000 477800 579400
rect 475200 577400 477800 578000
rect 475200 576000 475800 577400
rect 477200 576000 477800 577400
rect 475200 575400 477800 576000
rect 475200 574000 475800 575400
rect 477200 574000 477800 575400
rect 475200 573400 477800 574000
rect 475200 572000 475800 573400
rect 477200 572000 477800 573400
rect 475200 571400 477800 572000
rect 475200 570000 475800 571400
rect 477200 570000 477800 571400
rect 475200 569400 477800 570000
rect 475200 568000 475800 569400
rect 477200 568000 477800 569400
rect 475200 567400 477800 568000
rect 511690 574080 519090 574680
rect 511690 568680 512590 574080
rect 518490 568680 519090 574080
rect 511690 567980 519090 568680
rect 564280 574210 571680 574810
rect 564280 568810 565180 574210
rect 571080 568810 571680 574210
rect 564280 568110 571680 568810
rect 475200 566000 475800 567400
rect 477200 566000 477800 567400
rect 475200 565400 477800 566000
rect 475200 564000 475800 565400
rect 477200 564000 477800 565400
rect 475200 563400 477800 564000
rect 475200 562000 475800 563400
rect 477200 562000 477800 563400
rect 475200 561400 477800 562000
rect 475200 560000 475800 561400
rect 477200 560000 477800 561400
rect 475200 559400 477800 560000
rect 475200 558000 475800 559400
rect 477200 558000 477800 559400
rect 475200 557400 477800 558000
rect 475200 556000 475800 557400
rect 477200 556000 477800 557400
rect 475200 555400 477800 556000
rect 475200 554000 475800 555400
rect 477200 554000 477800 555400
rect 475200 553400 477800 554000
rect 475200 552000 475800 553400
rect 477200 552000 477800 553400
rect 475200 551400 477800 552000
rect 475200 550000 475800 551400
rect 477200 550000 477800 551400
rect 475200 549400 477800 550000
rect 475200 548000 475800 549400
rect 477200 548000 477800 549400
rect 475200 547400 477800 548000
rect 475200 546000 475800 547400
rect 477200 546000 477800 547400
rect 475200 545400 477800 546000
rect 475200 544400 475800 545400
rect 16800 544200 475800 544400
rect 15800 544000 475800 544200
rect 477200 544000 477800 545400
rect 511790 551080 519190 551780
rect 511790 545680 512790 551080
rect 518690 545680 519190 551080
rect 511790 545080 519190 545680
rect 564380 551210 571780 551910
rect 564380 545810 565380 551210
rect 571280 545810 571780 551210
rect 564380 545210 571780 545810
rect 15800 543400 477800 544000
rect 15800 542200 475800 543400
rect 15800 541800 17000 542200
rect 15800 541200 16000 541800
rect 16800 541200 17000 541800
rect 15800 538800 17000 541200
rect 15800 538200 16000 538800
rect 16800 538200 17000 538800
rect 3200 537600 5800 538000
rect 3200 536400 3800 537600
rect 5200 536400 5800 537600
rect 3200 535600 5800 536400
rect 3200 534400 3800 535600
rect 5200 534400 5800 535600
rect 3200 533600 5800 534400
rect 3200 532400 3800 533600
rect 5200 532400 5800 533600
rect 15800 535800 17000 538200
rect 15800 535200 16000 535800
rect 16800 535200 17000 535800
rect 10000 532800 10600 533200
rect 15800 532400 17000 535200
rect 475200 542000 475800 542200
rect 477200 542000 477800 543400
rect 475200 541400 477800 542000
rect 475200 540000 475800 541400
rect 477200 540000 477800 541400
rect 475200 539400 477800 540000
rect 475200 538000 475800 539400
rect 477200 538000 477800 539400
rect 475200 537400 477800 538000
rect 475200 536000 475800 537400
rect 477200 536000 477800 537400
rect 475200 535400 477800 536000
rect 475200 534000 475800 535400
rect 477200 534000 477800 535400
rect 475200 533400 477800 534000
rect 3200 531600 5800 532400
rect 3200 530400 3800 531600
rect 5200 530400 5800 531600
rect 3200 529600 5800 530400
rect 3200 528400 3800 529600
rect 5200 528400 5800 529600
rect 3200 527600 5800 528400
rect 10300 532200 17400 532400
rect 10300 531800 15800 532200
rect 17100 531800 17400 532200
rect 10300 531500 17400 531800
rect 10300 531100 15800 531500
rect 17100 531100 17400 531500
rect 10300 530900 17400 531100
rect 10300 530500 15800 530900
rect 17100 530500 17400 530900
rect 10300 530200 17400 530500
rect 10300 529800 15800 530200
rect 17100 529800 17400 530200
rect 10300 529500 17400 529800
rect 10300 529100 15800 529500
rect 17100 529100 17400 529500
rect 10300 528800 17400 529100
rect 10300 528400 15800 528800
rect 17100 528400 17400 528800
rect 10300 527800 17400 528400
rect 475200 532000 475800 533400
rect 477200 532000 477800 533400
rect 475200 531400 477800 532000
rect 491230 533850 499110 534220
rect 491230 532700 491350 533850
rect 499020 532700 499110 533850
rect 491230 531460 499110 532700
rect 543820 533980 551700 534350
rect 543820 532830 543940 533980
rect 551610 532830 551700 533980
rect 543820 531590 551700 532830
rect 475200 530000 475800 531400
rect 477200 530000 477800 531400
rect 475200 529400 477800 530000
rect 475200 528000 475800 529400
rect 477200 528000 477800 529400
rect 3200 526400 3800 527600
rect 5200 526400 5800 527600
rect 10000 527000 10600 527400
rect 15800 527200 17000 527800
rect 3200 525600 5800 526400
rect 3200 524400 3800 525600
rect 5200 524400 5800 525600
rect 3200 523600 5800 524400
rect 3200 522400 3800 523600
rect 5200 522400 5800 523600
rect 3200 521600 5800 522400
rect 3200 520400 3800 521600
rect 5200 520400 5800 521600
rect 3200 519600 5800 520400
rect 3200 518400 3800 519600
rect 5200 518400 5800 519600
rect 3200 517600 5800 518400
rect 3200 516400 3800 517600
rect 5200 516400 5800 517600
rect 3200 515600 5800 516400
rect 3200 514400 3800 515600
rect 5200 514400 5800 515600
rect 3200 513600 5800 514400
rect 3200 512400 3800 513600
rect 5200 512400 5800 513600
rect 3200 511600 5800 512400
rect 3200 510400 3800 511600
rect 5200 510400 5800 511600
rect 3200 509600 5800 510400
rect 3200 508400 3800 509600
rect 5200 508400 5800 509600
rect 3200 507600 5800 508400
rect 3200 506400 3800 507600
rect 5200 506400 5800 507600
rect 3200 505600 5800 506400
rect 3200 504400 3800 505600
rect 5200 504400 5800 505600
rect 3200 503600 5800 504400
rect 3200 502400 3800 503600
rect 5200 502400 5800 503600
rect 3200 501600 5800 502400
rect 3200 500400 3800 501600
rect 5200 500400 5800 501600
rect 3200 499600 5800 500400
rect 3200 498400 3800 499600
rect 5200 498400 5800 499600
rect 3200 497600 5800 498400
rect 3200 496400 3800 497600
rect 5200 496400 5800 497600
rect 3200 495600 5800 496400
rect 3200 494400 3800 495600
rect 5200 494400 5800 495600
rect 3200 493600 5800 494400
rect 3200 492400 3800 493600
rect 5200 492400 5800 493600
rect 3200 491600 5800 492400
rect 3200 490400 3800 491600
rect 5200 490400 5800 491600
rect 3200 489600 5800 490400
rect 3200 488400 3800 489600
rect 5200 488400 5800 489600
rect 3200 487600 5800 488400
rect 3200 486400 3800 487600
rect 5200 486400 5800 487600
rect 3200 485600 5800 486400
rect 3200 484400 3800 485600
rect 5200 484400 5800 485600
rect 3200 483600 5800 484400
rect 3200 482400 3800 483600
rect 5200 482400 5800 483600
rect 3200 481600 5800 482400
rect 3200 480400 3800 481600
rect 5200 480400 5800 481600
rect 3200 479600 5800 480400
rect 3200 478400 3800 479600
rect 5200 478400 5800 479600
rect 3200 477600 5800 478400
rect 3200 476400 3800 477600
rect 5200 476400 5800 477600
rect 3200 475600 5800 476400
rect 3200 474400 3800 475600
rect 5200 474400 5800 475600
rect 3200 473600 5800 474400
rect 3200 472400 3800 473600
rect 5200 472400 5800 473600
rect 3200 471600 5800 472400
rect 3200 470400 3800 471600
rect 5200 470400 5800 471600
rect 3200 469600 5800 470400
rect 3200 468400 3800 469600
rect 5200 468400 5800 469600
rect 3200 467600 5800 468400
rect 3200 466400 3800 467600
rect 5200 466400 5800 467600
rect 3200 465600 5800 466400
rect 3200 464400 3800 465600
rect 5200 464400 5800 465600
rect 3200 463600 5800 464400
rect 3200 462400 3800 463600
rect 5200 462400 5800 463600
rect 3200 461600 5800 462400
rect 3200 460400 3800 461600
rect 5200 460400 5800 461600
rect 3200 459600 5800 460400
rect 3200 458400 3800 459600
rect 5200 458400 5800 459600
rect 3200 457600 5800 458400
rect 3200 456400 3800 457600
rect 5200 456400 5800 457600
rect 3200 455600 5800 456400
rect 3200 454400 3800 455600
rect 5200 454400 5800 455600
rect 3200 453600 5800 454400
rect 3200 452400 3800 453600
rect 5200 452400 5800 453600
rect 3200 451600 5800 452400
rect 3200 450400 3800 451600
rect 5200 450400 5800 451600
rect 3200 449600 5800 450400
rect 3200 448400 3800 449600
rect 5200 448400 5800 449600
rect 3200 447600 5800 448400
rect 3200 446400 3800 447600
rect 5200 446400 5800 447600
rect 3200 445600 5800 446400
rect 3200 444400 3800 445600
rect 5200 444400 5800 445600
rect 3200 443600 5800 444400
rect 3200 442400 3800 443600
rect 5200 442400 5800 443600
rect 3200 441600 5800 442400
rect 3200 440400 3800 441600
rect 5200 440400 5800 441600
rect 3200 439600 5800 440400
rect 3200 438400 3800 439600
rect 5200 438400 5800 439600
rect 3200 437600 5800 438400
rect 3200 436400 3800 437600
rect 5200 436400 5800 437600
rect 3200 435600 5800 436400
rect 3200 434400 3800 435600
rect 5200 434400 5800 435600
rect 3200 433600 5800 434400
rect 3200 432400 3800 433600
rect 5200 432400 5800 433600
rect 3200 375600 5800 432400
rect 600 375400 5800 375600
rect 600 375000 1000 375400
rect 2000 375000 5800 375400
rect 600 374800 5800 375000
rect 600 374400 1000 374800
rect 2000 374400 5800 374800
rect 600 374000 5800 374400
rect 600 373600 1000 374000
rect 2000 373600 5800 374000
rect 600 373200 5800 373600
rect 600 372800 1000 373200
rect 2000 372800 5800 373200
rect 600 372400 5800 372800
rect 600 372000 1000 372400
rect 2000 372000 5800 372400
rect 600 371600 5800 372000
rect 600 371200 1000 371600
rect 2000 371200 5800 371600
rect 600 370800 5800 371200
rect 600 370400 1000 370800
rect 2000 370400 5800 370800
rect 600 370000 5800 370400
rect 15800 526600 16000 527200
rect 16800 526600 17000 527200
rect 15800 524200 17000 526600
rect 15800 523600 16000 524200
rect 16800 523600 17000 524200
rect 15800 521200 17000 523600
rect 15800 520600 16000 521200
rect 16800 520600 17000 521200
rect 15800 518200 17000 520600
rect 15800 517600 16000 518200
rect 16800 517600 17000 518200
rect 15800 515200 17000 517600
rect 15800 514600 16000 515200
rect 16800 514600 17000 515200
rect 15800 512200 17000 514600
rect 15800 511600 16000 512200
rect 16800 511600 17000 512200
rect 15800 509200 17000 511600
rect 15800 508600 16000 509200
rect 16800 508600 17000 509200
rect 15800 506200 17000 508600
rect 15800 505600 16000 506200
rect 16800 505600 17000 506200
rect 15800 503200 17000 505600
rect 15800 502600 16000 503200
rect 16800 502600 17000 503200
rect 15800 500200 17000 502600
rect 15800 499600 16000 500200
rect 16800 499600 17000 500200
rect 15800 497200 17000 499600
rect 15800 496600 16000 497200
rect 16800 496600 17000 497200
rect 15800 494200 17000 496600
rect 15800 493600 16000 494200
rect 16800 493600 17000 494200
rect 15800 491200 17000 493600
rect 15800 490600 16000 491200
rect 16800 490600 17000 491200
rect 15800 488200 17000 490600
rect 15800 487600 16000 488200
rect 16800 487600 17000 488200
rect 15800 485200 17000 487600
rect 15800 484600 16000 485200
rect 16800 484600 17000 485200
rect 15800 482200 17000 484600
rect 15800 481600 16000 482200
rect 16800 481600 17000 482200
rect 15800 479200 17000 481600
rect 15800 478600 16000 479200
rect 16800 478600 17000 479200
rect 15800 476200 17000 478600
rect 15800 475600 16000 476200
rect 16800 475600 17000 476200
rect 15800 473200 17000 475600
rect 15800 472600 16000 473200
rect 16800 472600 17000 473200
rect 15800 470200 17000 472600
rect 15800 469600 16000 470200
rect 16800 469600 17000 470200
rect 15800 467200 17000 469600
rect 15800 466600 16000 467200
rect 16800 466600 17000 467200
rect 15800 464200 17000 466600
rect 15800 463600 16000 464200
rect 16800 463600 17000 464200
rect 15800 461200 17000 463600
rect 15800 460600 16000 461200
rect 16800 460600 17000 461200
rect 15800 458200 17000 460600
rect 15800 457600 16000 458200
rect 16800 457600 17000 458200
rect 15800 455200 17000 457600
rect 15800 454600 16000 455200
rect 16800 454600 17000 455200
rect 15800 452200 17000 454600
rect 15800 451600 16000 452200
rect 16800 451600 17000 452200
rect 15800 449200 17000 451600
rect 15800 448600 16000 449200
rect 16800 448600 17000 449200
rect 15800 446200 17000 448600
rect 15800 445600 16000 446200
rect 16800 445600 17000 446200
rect 15800 443200 17000 445600
rect 15800 442600 16000 443200
rect 16800 442600 17000 443200
rect 15800 440200 17000 442600
rect 15800 439600 16000 440200
rect 16800 439600 17000 440200
rect 15800 437200 17000 439600
rect 15800 436600 16000 437200
rect 16800 436600 17000 437200
rect 15800 434200 17000 436600
rect 15800 433600 16000 434200
rect 16800 433600 17000 434200
rect 15800 431200 17000 433600
rect 15800 430600 16000 431200
rect 16800 430600 17000 431200
rect 15800 428200 17000 430600
rect 15800 427600 16000 428200
rect 16800 427600 17000 428200
rect 15800 425200 17000 427600
rect 15800 424600 16000 425200
rect 16800 424600 17000 425200
rect 15800 422200 17000 424600
rect 15800 421600 16000 422200
rect 16800 421600 17000 422200
rect 15800 419200 17000 421600
rect 15800 418600 16000 419200
rect 16800 418600 17000 419200
rect 15800 416200 17000 418600
rect 15800 415600 16000 416200
rect 16800 415600 17000 416200
rect 15800 413200 17000 415600
rect 15800 412600 16000 413200
rect 16800 412600 17000 413200
rect 15800 410200 17000 412600
rect 15800 409600 16000 410200
rect 16800 409600 17000 410200
rect 15800 407200 17000 409600
rect 15800 406600 16000 407200
rect 16800 406600 17000 407200
rect 15800 404200 17000 406600
rect 15800 403600 16000 404200
rect 16800 403600 17000 404200
rect 15800 401200 17000 403600
rect 15800 400600 16000 401200
rect 16800 400600 17000 401200
rect 15800 398200 17000 400600
rect 15800 397600 16000 398200
rect 16800 397600 17000 398200
rect 15800 395200 17000 397600
rect 15800 394600 16000 395200
rect 16800 394600 17000 395200
rect 15800 392200 17000 394600
rect 15800 391600 16000 392200
rect 16800 391600 17000 392200
rect 15800 389200 17000 391600
rect 15800 388600 16000 389200
rect 16800 388600 17000 389200
rect 15800 386200 17000 388600
rect 15800 385600 16000 386200
rect 16800 385600 17000 386200
rect 15800 383200 17000 385600
rect 15800 382600 16000 383200
rect 16800 382600 17000 383200
rect 15800 380200 17000 382600
rect 15800 379600 16000 380200
rect 16800 379600 17000 380200
rect 15800 377200 17000 379600
rect 15800 376600 16000 377200
rect 16800 376600 17000 377200
rect 15800 374200 17000 376600
rect 15800 373600 16000 374200
rect 16800 373600 17000 374200
rect 15800 371200 17000 373600
rect 15800 370600 16000 371200
rect 16800 370600 17000 371200
rect 600 369400 1600 370000
rect 600 368800 800 369400
rect 1400 368800 1600 369400
rect 600 367400 1600 368800
rect 600 366800 800 367400
rect 1400 366800 1600 367400
rect 600 365400 1600 366800
rect 600 364800 800 365400
rect 1400 364800 1600 365400
rect 600 363400 1600 364800
rect 600 362800 800 363400
rect 1400 362800 1600 363400
rect 600 361400 1600 362800
rect 600 360800 800 361400
rect 1400 360800 1600 361400
rect 600 359400 1600 360800
rect 600 358800 800 359400
rect 1400 358800 1600 359400
rect 600 357400 1600 358800
rect 600 356800 800 357400
rect 1400 356800 1600 357400
rect 600 355400 1600 356800
rect 600 354800 800 355400
rect 1400 354800 1600 355400
rect 600 353400 1600 354800
rect 600 352800 800 353400
rect 1400 352800 1600 353400
rect 600 351400 1600 352800
rect 600 350800 800 351400
rect 1400 350800 1600 351400
rect 600 349400 1600 350800
rect 600 348800 800 349400
rect 1400 348800 1600 349400
rect 600 347400 1600 348800
rect 600 346800 800 347400
rect 1400 346800 1600 347400
rect 600 345400 1600 346800
rect 600 344800 800 345400
rect 1400 344800 1600 345400
rect 600 344200 1600 344800
rect 15800 341800 17000 370600
rect 15800 341200 16000 341800
rect 16800 341200 17000 341800
rect 13800 339300 14143 339600
rect 15800 338800 17000 341200
rect 13800 338300 14143 338600
rect 15800 338200 16000 338800
rect 16800 338200 17000 338800
rect 13800 337300 14143 337600
rect 13800 336300 14143 336600
rect 15800 335800 17000 338200
rect 13800 335300 14143 335600
rect 15800 335200 16000 335800
rect 16800 335200 17000 335800
rect 13800 334300 14143 334600
rect 13800 333300 14143 333600
rect 15800 332800 17000 335200
rect 15800 332200 16000 332800
rect 16800 332200 17000 332800
rect 15800 329800 17000 332200
rect 15800 329200 16000 329800
rect 16800 329200 17000 329800
rect 15800 326800 17000 329200
rect 15800 326200 16000 326800
rect 16800 326200 17000 326800
rect 15800 323800 17000 326200
rect 15800 323200 16000 323800
rect 16800 323200 17000 323800
rect 15800 320800 17000 323200
rect 15800 320200 16000 320800
rect 16800 320200 17000 320800
rect 15800 317800 17000 320200
rect 15800 317200 16000 317800
rect 16800 317200 17000 317800
rect 15800 314800 17000 317200
rect 15800 314200 16000 314800
rect 16800 314200 17000 314800
rect 15800 311800 17000 314200
rect 15800 311200 16000 311800
rect 16800 311200 17000 311800
rect 15800 308800 17000 311200
rect 15800 308200 16000 308800
rect 16800 308200 17000 308800
rect 15800 305800 17000 308200
rect 15800 305200 16000 305800
rect 16800 305200 17000 305800
rect 15800 302800 17000 305200
rect 15800 302200 16000 302800
rect 16800 302200 17000 302800
rect 15800 299800 17000 302200
rect 15800 299200 16000 299800
rect 16800 299200 17000 299800
rect 15800 296800 17000 299200
rect 15800 296200 16000 296800
rect 16800 296200 17000 296800
rect 15800 293800 17000 296200
rect 15800 293200 16000 293800
rect 16800 293200 17000 293800
rect 15800 290800 17000 293200
rect 15800 290200 16000 290800
rect 16800 290200 17000 290800
rect 15800 287800 17000 290200
rect 15800 287200 16000 287800
rect 16800 287200 17000 287800
rect 15800 284800 17000 287200
rect 15800 284200 16000 284800
rect 16800 284200 17000 284800
rect 15800 281800 17000 284200
rect 15800 281200 16000 281800
rect 16800 281200 17000 281800
rect 15800 278800 17000 281200
rect 15800 278200 16000 278800
rect 16800 278200 17000 278800
rect 15800 275800 17000 278200
rect 15800 275200 16000 275800
rect 16800 275200 17000 275800
rect 15800 272800 17000 275200
rect 15800 272200 16000 272800
rect 16800 272200 17000 272800
rect 15800 269800 17000 272200
rect 15800 269200 16000 269800
rect 16800 269200 17000 269800
rect 15800 266800 17000 269200
rect 15800 266200 16000 266800
rect 16800 266200 17000 266800
rect 15800 263800 17000 266200
rect 15800 263200 16000 263800
rect 16800 263200 17000 263800
rect 15800 260800 17000 263200
rect 15800 260200 16000 260800
rect 16800 260200 17000 260800
rect 15800 257800 17000 260200
rect 15800 257200 16000 257800
rect 16800 257200 17000 257800
rect 15800 254800 17000 257200
rect 15800 254200 16000 254800
rect 16800 254200 17000 254800
rect 15800 251800 17000 254200
rect 15800 251200 16000 251800
rect 16800 251200 17000 251800
rect 15800 248800 17000 251200
rect 15800 248200 16000 248800
rect 16800 248200 17000 248800
rect 15800 245800 17000 248200
rect 15800 245200 16000 245800
rect 16800 245200 17000 245800
rect 15800 242800 17000 245200
rect 15800 242200 16000 242800
rect 16800 242200 17000 242800
rect 15800 239800 17000 242200
rect 15800 239200 16000 239800
rect 16800 239200 17000 239800
rect 15800 236800 17000 239200
rect 15800 236200 16000 236800
rect 16800 236200 17000 236800
rect 15800 233800 17000 236200
rect 15800 233200 16000 233800
rect 16800 233200 17000 233800
rect 15800 230800 17000 233200
rect 15800 230200 16000 230800
rect 16800 230200 17000 230800
rect 15800 227800 17000 230200
rect 15800 227200 16000 227800
rect 16800 227200 17000 227800
rect 15800 224800 17000 227200
rect 15800 224200 16000 224800
rect 16800 224200 17000 224800
rect 15800 221800 17000 224200
rect 15800 221200 16000 221800
rect 16800 221200 17000 221800
rect 15800 218800 17000 221200
rect 15800 218200 16000 218800
rect 16800 218200 17000 218800
rect 15800 215800 17000 218200
rect 15800 215200 16000 215800
rect 16800 215200 17000 215800
rect 15800 212800 17000 215200
rect 15800 212200 16000 212800
rect 16800 212200 17000 212800
rect 15800 209800 17000 212200
rect 15800 209200 16000 209800
rect 16800 209200 17000 209800
rect 15800 206800 17000 209200
rect 15800 206200 16000 206800
rect 16800 206200 17000 206800
rect 15800 203800 17000 206200
rect 15800 203200 16000 203800
rect 16800 203200 17000 203800
rect 15800 200800 17000 203200
rect 15800 200200 16000 200800
rect 16800 200200 17000 200800
rect 15800 197800 17000 200200
rect 15800 197200 16000 197800
rect 16800 197200 17000 197800
rect 15800 194800 17000 197200
rect 15800 194200 16000 194800
rect 16800 194200 17000 194800
rect 15800 191800 17000 194200
rect 15800 191200 16000 191800
rect 16800 191200 17000 191800
rect 15800 188800 17000 191200
rect 15800 188200 16000 188800
rect 16800 188200 17000 188800
rect 15800 185800 17000 188200
rect 15800 185200 16000 185800
rect 16800 185200 17000 185800
rect 15800 182800 17000 185200
rect 15800 182200 16000 182800
rect 16800 182200 17000 182800
rect 15800 179800 17000 182200
rect 15800 179200 16000 179800
rect 16800 179200 17000 179800
rect 400 177370 2740 177720
rect 400 163110 700 177370
rect 2330 163110 2740 177370
rect 400 162870 2740 163110
rect 15800 176800 17000 179200
rect 15800 176200 16000 176800
rect 16800 176200 17000 176800
rect 15800 173800 17000 176200
rect 15800 173200 16000 173800
rect 16800 173200 17000 173800
rect 15800 170800 17000 173200
rect 15800 170200 16000 170800
rect 16800 170200 17000 170800
rect 15800 167800 17000 170200
rect 15800 167200 16000 167800
rect 16800 167200 17000 167800
rect 15800 164800 17000 167200
rect 15800 164200 16000 164800
rect 16800 164200 17000 164800
rect 15800 161800 17000 164200
rect 15800 161200 16000 161800
rect 16800 161200 17000 161800
rect 15800 158800 17000 161200
rect 15800 158200 16000 158800
rect 16800 158200 17000 158800
rect 15800 155800 17000 158200
rect 15800 155200 16000 155800
rect 16800 155200 17000 155800
rect 15800 152800 17000 155200
rect 15800 152200 16000 152800
rect 16800 152200 17000 152800
rect 15800 149800 17000 152200
rect 15800 149200 16000 149800
rect 16800 149200 17000 149800
rect 15800 146800 17000 149200
rect 15800 146200 16000 146800
rect 16800 146200 17000 146800
rect 15800 143800 17000 146200
rect 15800 143200 16000 143800
rect 16800 143200 17000 143800
rect 15800 140800 17000 143200
rect 15800 140200 16000 140800
rect 16800 140200 17000 140800
rect 15800 137800 17000 140200
rect 15800 137200 16000 137800
rect 16800 137200 17000 137800
rect 15800 134800 17000 137200
rect 15800 134200 16000 134800
rect 16800 134200 17000 134800
rect 15800 131800 17000 134200
rect 15800 131200 16000 131800
rect 16800 131200 17000 131800
rect 15800 128800 17000 131200
rect 15800 128200 16000 128800
rect 16800 128200 17000 128800
rect 15800 125800 17000 128200
rect 15800 125200 16000 125800
rect 16800 125200 17000 125800
rect 15800 122800 17000 125200
rect 15800 122200 16000 122800
rect 16800 122200 17000 122800
rect 15800 119800 17000 122200
rect 15800 119200 16000 119800
rect 16800 119200 17000 119800
rect 15800 116800 17000 119200
rect 15800 116200 16000 116800
rect 16800 116200 17000 116800
rect 15800 113800 17000 116200
rect 15800 113200 16000 113800
rect 16800 113200 17000 113800
rect 15800 110800 17000 113200
rect 15800 110200 16000 110800
rect 16800 110200 17000 110800
rect 15800 107800 17000 110200
rect 15800 107200 16000 107800
rect 16800 107200 17000 107800
rect 15800 104800 17000 107200
rect 15800 104200 16000 104800
rect 16800 104200 17000 104800
rect 15800 101800 17000 104200
rect 15800 101200 16000 101800
rect 16800 101200 17000 101800
rect 15800 98800 17000 101200
rect 15800 98200 16000 98800
rect 16800 98200 17000 98800
rect 15800 95800 17000 98200
rect 15800 95200 16000 95800
rect 16800 95200 17000 95800
rect 15800 92800 17000 95200
rect 15800 92200 16000 92800
rect 16800 92200 17000 92800
rect 15800 89800 17000 92200
rect 15800 89200 16000 89800
rect 16800 89200 17000 89800
rect 15800 86800 17000 89200
rect 15800 86200 16000 86800
rect 16800 86200 17000 86800
rect 15800 83800 17000 86200
rect 15800 83200 16000 83800
rect 16800 83200 17000 83800
rect 15800 80800 17000 83200
rect 15800 80200 16000 80800
rect 16800 80200 17000 80800
rect 15800 77800 17000 80200
rect 15800 77200 16000 77800
rect 16800 77200 17000 77800
rect 15800 74800 17000 77200
rect 15800 74200 16000 74800
rect 16800 74200 17000 74800
rect 15800 71800 17000 74200
rect 15800 71200 16000 71800
rect 16800 71200 17000 71800
rect 15800 68800 17000 71200
rect 15800 68200 16000 68800
rect 16800 68200 17000 68800
rect 15800 65800 17000 68200
rect 15800 65200 16000 65800
rect 16800 65200 17000 65800
rect 15800 62800 17000 65200
rect 15800 62200 16000 62800
rect 16800 62200 17000 62800
rect 15800 59800 17000 62200
rect 15800 59200 16000 59800
rect 16800 59200 17000 59800
rect 15800 56800 17000 59200
rect 15800 56200 16000 56800
rect 16800 56200 17000 56800
rect 15800 53800 17000 56200
rect 15800 53200 16000 53800
rect 16800 53200 17000 53800
rect 15800 50800 17000 53200
rect 15800 50200 16000 50800
rect 16800 50200 17000 50800
rect 15800 47800 17000 50200
rect 15800 47200 16000 47800
rect 16800 47200 17000 47800
rect 15800 44800 17000 47200
rect 15800 44200 16000 44800
rect 16800 44200 17000 44800
rect 15800 41800 17000 44200
rect 15800 41200 16000 41800
rect 16800 41200 17000 41800
rect 15800 38800 17000 41200
rect 15800 38200 16000 38800
rect 16800 38200 17000 38800
rect 15800 35800 17000 38200
rect 15800 35200 16000 35800
rect 16800 35200 17000 35800
rect 15800 32800 17000 35200
rect 15800 32200 16000 32800
rect 16800 32200 17000 32800
rect 15800 29800 17000 32200
rect 15800 29200 16000 29800
rect 16800 29200 17000 29800
rect 15800 26800 17000 29200
rect 15800 26200 16000 26800
rect 16800 26200 17000 26800
rect 15800 23800 17000 26200
rect 15800 23200 16000 23800
rect 16800 23200 17000 23800
rect 15800 20800 17000 23200
rect 15800 20200 16000 20800
rect 16800 20200 17000 20800
rect 15800 17800 17000 20200
rect 15800 17200 16000 17800
rect 16800 17200 17000 17800
rect 15800 14800 17000 17200
rect 15800 14200 16000 14800
rect 16800 14200 17000 14800
rect 15800 11800 17000 14200
rect 15800 11200 16000 11800
rect 16800 11200 17000 11800
rect 15800 8800 17000 11200
rect 15800 8200 16000 8800
rect 16800 8200 17000 8800
rect 15800 5800 17000 8200
rect 15800 5200 16000 5800
rect 16800 5200 17000 5800
rect 15800 4400 17000 5200
rect 475200 527400 477800 528000
rect 475200 526000 475800 527400
rect 477200 526000 477800 527400
rect 475200 525400 477800 526000
rect 475200 524000 475800 525400
rect 477200 524000 477800 525400
rect 475200 523400 477800 524000
rect 475200 522000 475800 523400
rect 477200 522000 477800 523400
rect 475200 521400 477800 522000
rect 475200 520000 475800 521400
rect 477200 520000 477800 521400
rect 511890 527380 519190 528080
rect 511890 522080 512590 527380
rect 518590 522080 519190 527380
rect 511890 521380 519190 522080
rect 564480 527510 571780 528210
rect 564480 522210 565180 527510
rect 571180 522210 571780 527510
rect 564480 521510 571780 522210
rect 475200 519400 477800 520000
rect 475200 518000 475800 519400
rect 477200 518000 477800 519400
rect 475200 517400 477800 518000
rect 475200 516000 475800 517400
rect 477200 516000 477800 517400
rect 475200 515400 477800 516000
rect 475200 514000 475800 515400
rect 477200 514000 477800 515400
rect 475200 513400 477800 514000
rect 475200 512000 475800 513400
rect 477200 512000 477800 513400
rect 475200 511400 477800 512000
rect 475200 510000 475800 511400
rect 477200 510000 477800 511400
rect 475200 509400 477800 510000
rect 475200 508000 475800 509400
rect 477200 508000 477800 509400
rect 475200 507400 477800 508000
rect 475200 506000 475800 507400
rect 477200 506000 477800 507400
rect 475200 505400 477800 506000
rect 475200 504000 475800 505400
rect 477200 504000 477800 505400
rect 475200 503400 477800 504000
rect 475200 502000 475800 503400
rect 477200 502000 477800 503400
rect 475200 501400 477800 502000
rect 475200 500000 475800 501400
rect 477200 500000 477800 501400
rect 475200 499400 477800 500000
rect 475200 498000 475800 499400
rect 477200 498000 477800 499400
rect 475200 497400 477800 498000
rect 475200 496000 475800 497400
rect 477200 496000 477800 497400
rect 475200 495400 477800 496000
rect 475200 494000 475800 495400
rect 477200 494000 477800 495400
rect 475200 493400 477800 494000
rect 475200 492000 475800 493400
rect 477200 492000 477800 493400
rect 528170 500750 530930 500870
rect 528170 493080 529410 500750
rect 530560 493080 530930 500750
rect 528170 492990 530930 493080
rect 475200 491400 477800 492000
rect 475200 490000 475800 491400
rect 477200 490000 477800 491400
rect 475200 489400 477800 490000
rect 475200 488000 475800 489400
rect 477200 488000 477800 489400
rect 475200 487400 477800 488000
rect 475200 486000 475800 487400
rect 477200 486000 477800 487400
rect 475200 485400 477800 486000
rect 475200 484000 475800 485400
rect 477200 484000 477800 485400
rect 475200 483400 477800 484000
rect 475200 482000 475800 483400
rect 477200 482000 477800 483400
rect 475200 481400 477800 482000
rect 475200 480000 475800 481400
rect 477200 480000 477800 481400
rect 475200 479400 477800 480000
rect 475200 478000 475800 479400
rect 477200 478000 477800 479400
rect 475200 477400 477800 478000
rect 475200 476000 475800 477400
rect 477200 476000 477800 477400
rect 475200 475400 477800 476000
rect 475200 474000 475800 475400
rect 477200 474000 477800 475400
rect 475200 473400 477800 474000
rect 475200 472000 475800 473400
rect 477200 472000 477800 473400
rect 518090 479510 524790 480210
rect 518090 473510 518790 479510
rect 524090 473510 524790 479510
rect 518090 472910 524790 473510
rect 541790 479310 548490 480310
rect 541790 473410 542390 479310
rect 547790 473410 548490 479310
rect 541790 472910 548490 473410
rect 564690 479510 571390 480410
rect 564690 473610 565390 479510
rect 570790 473610 571390 479510
rect 564690 473010 571390 473610
rect 475200 471400 477800 472000
rect 475200 470000 475800 471400
rect 477200 470000 477800 471400
rect 475200 469400 477800 470000
rect 475200 468000 475800 469400
rect 477200 468000 477800 469400
rect 475200 467400 477800 468000
rect 475200 466000 475800 467400
rect 477200 466000 477800 467400
rect 475200 465400 477800 466000
rect 475200 464000 475800 465400
rect 477200 464000 477800 465400
rect 475200 463400 477800 464000
rect 475200 462000 475800 463400
rect 477200 463000 477800 463400
rect 477200 462000 478600 463000
rect 475200 461400 478600 462000
rect 475200 460000 475800 461400
rect 477200 460000 478600 461400
rect 475200 459400 478600 460000
rect 475200 458000 475800 459400
rect 477200 458000 478600 459400
rect 475200 457400 478600 458000
rect 475200 456000 475800 457400
rect 477200 456000 478600 457400
rect 475200 455400 478600 456000
rect 475200 454000 475800 455400
rect 477200 454000 478600 455400
rect 475200 453400 478600 454000
rect 475200 452000 475800 453400
rect 477200 452000 478600 453400
rect 475200 451400 478600 452000
rect 475200 450000 475800 451400
rect 477200 450000 478600 451400
rect 475200 449400 478600 450000
rect 475200 448000 475800 449400
rect 477200 448000 478600 449400
rect 475200 447400 478600 448000
rect 475200 446000 475800 447400
rect 477200 446000 478600 447400
rect 475200 445400 478600 446000
rect 475200 444000 475800 445400
rect 477200 444000 478600 445400
rect 475200 443400 478600 444000
rect 475200 442000 475800 443400
rect 477200 442000 478600 443400
rect 475200 441400 478600 442000
rect 475200 440000 475800 441400
rect 477200 440000 478600 441400
rect 475200 439400 478600 440000
rect 475200 438000 475800 439400
rect 477200 438000 478600 439400
rect 475200 437400 478600 438000
rect 475200 436000 475800 437400
rect 477200 436000 478600 437400
rect 475200 435400 478600 436000
rect 475200 434000 475800 435400
rect 477200 434000 478600 435400
rect 475200 433400 478600 434000
rect 475200 432000 475800 433400
rect 477200 432000 478600 433400
rect 475200 431400 478600 432000
rect 475200 430000 475800 431400
rect 477200 430000 478600 431400
rect 475200 429400 478600 430000
rect 475200 428000 475800 429400
rect 477200 428000 478600 429400
rect 475200 427400 478600 428000
rect 475200 426000 475800 427400
rect 477200 426000 478600 427400
rect 475200 425400 478600 426000
rect 475200 424000 475800 425400
rect 477200 424000 478600 425400
rect 475200 423400 478600 424000
rect 475200 422000 475800 423400
rect 477200 422000 478600 423400
rect 475200 421400 478600 422000
rect 475200 420000 475800 421400
rect 477200 420000 478600 421400
rect 475200 419400 478600 420000
rect 475200 418000 475800 419400
rect 477200 418000 478600 419400
rect 475200 417400 478600 418000
rect 475200 416000 475800 417400
rect 477200 416000 478600 417400
rect 475200 415400 478600 416000
rect 475200 414000 475800 415400
rect 477200 414000 478600 415400
rect 475200 413400 478600 414000
rect 475200 412000 475800 413400
rect 477200 412000 478600 413400
rect 475200 411400 478600 412000
rect 475200 410000 475800 411400
rect 477200 410000 478600 411400
rect 475200 409400 478600 410000
rect 475200 408000 475800 409400
rect 477200 408000 478600 409400
rect 475200 407400 478600 408000
rect 475200 406000 475800 407400
rect 477200 406000 478600 407400
rect 475200 405400 478600 406000
rect 475200 404000 475800 405400
rect 477200 404000 478600 405400
rect 475200 403400 478600 404000
rect 475200 402000 475800 403400
rect 477200 402000 478600 403400
rect 475200 401400 478600 402000
rect 475200 400000 475800 401400
rect 477200 400000 478600 401400
rect 475200 399400 478600 400000
rect 475200 398000 475800 399400
rect 477200 398000 478600 399400
rect 475200 397400 478600 398000
rect 475200 396000 475800 397400
rect 477200 396000 478600 397400
rect 475200 395400 478600 396000
rect 475200 394000 475800 395400
rect 477200 394000 478600 395400
rect 475200 393400 478600 394000
rect 475200 392000 475800 393400
rect 477200 392000 478600 393400
rect 475200 391400 478600 392000
rect 475200 390000 475800 391400
rect 477200 390000 478600 391400
rect 475200 389400 478600 390000
rect 475200 388000 475800 389400
rect 477200 388000 478600 389400
rect 475200 387400 478600 388000
rect 475200 386000 475800 387400
rect 477200 386000 478600 387400
rect 475200 385400 478600 386000
rect 475200 384000 475800 385400
rect 477200 384000 478600 385400
rect 475200 383400 478600 384000
rect 475200 382000 475800 383400
rect 477200 382000 478600 383400
rect 475200 381400 478600 382000
rect 475200 380000 475800 381400
rect 477200 380000 478600 381400
rect 475200 379400 478600 380000
rect 475200 378000 475800 379400
rect 477200 378000 478600 379400
rect 475200 377400 478600 378000
rect 475200 376000 475800 377400
rect 477200 376000 478600 377400
rect 475200 375400 478600 376000
rect 475200 374000 475800 375400
rect 477200 374000 478600 375400
rect 475200 373400 478600 374000
rect 475200 372000 475800 373400
rect 477200 372400 478600 373400
rect 576400 396400 582600 397600
rect 576400 395800 576800 396400
rect 582200 395800 582600 396400
rect 576400 394400 582600 395800
rect 576400 393800 576800 394400
rect 582200 393800 582600 394400
rect 576400 392400 582600 393800
rect 576400 391800 576800 392400
rect 582200 391800 582600 392400
rect 576400 390400 582600 391800
rect 576400 389800 576800 390400
rect 582200 389800 582600 390400
rect 576400 388400 582600 389800
rect 576400 387800 576800 388400
rect 582200 387800 582600 388400
rect 576400 386400 582600 387800
rect 576400 385800 576800 386400
rect 582200 385800 582600 386400
rect 576400 384400 582600 385800
rect 576400 383800 576800 384400
rect 582200 383800 582600 384400
rect 576400 382400 582600 383800
rect 576400 381800 576800 382400
rect 582200 381800 582600 382400
rect 576400 380400 582600 381800
rect 576400 379800 576800 380400
rect 582200 379800 582600 380400
rect 576400 378400 582600 379800
rect 576400 377800 576800 378400
rect 582200 377800 582600 378400
rect 576400 376400 582600 377800
rect 576400 375800 576800 376400
rect 582200 375800 582600 376400
rect 576400 374400 582600 375800
rect 576400 373800 576800 374400
rect 582200 373800 582600 374400
rect 576400 372400 582600 373800
rect 477200 372000 576800 372400
rect 475200 371800 576800 372000
rect 582200 371800 582600 372400
rect 475200 371400 582600 371800
rect 475200 370000 475800 371400
rect 477200 370400 582600 371400
rect 477200 370000 576800 370400
rect 475200 369800 576800 370000
rect 582200 369800 582600 370400
rect 475200 369400 582600 369800
rect 475200 368000 475800 369400
rect 477200 368000 478600 369400
rect 475200 367400 478600 368000
rect 475200 366000 475800 367400
rect 477200 366000 478600 367400
rect 475200 365400 478600 366000
rect 475200 364000 475800 365400
rect 477200 364000 478600 365400
rect 475200 363400 478600 364000
rect 475200 362000 475800 363400
rect 477200 362000 478600 363400
rect 475200 361400 478600 362000
rect 475200 360000 475800 361400
rect 477200 360000 478600 361400
rect 475200 359400 478600 360000
rect 475200 358000 475800 359400
rect 477200 358000 478600 359400
rect 475200 357400 478600 358000
rect 475200 356000 475800 357400
rect 477200 356000 478600 357400
rect 475200 355400 478600 356000
rect 475200 354000 475800 355400
rect 477200 354000 478600 355400
rect 475200 353400 478600 354000
rect 475200 352000 475800 353400
rect 477200 352000 478600 353400
rect 475200 351400 478600 352000
rect 475200 350000 475800 351400
rect 477200 350000 478600 351400
rect 475200 349400 478600 350000
rect 475200 348000 475800 349400
rect 477200 348000 478600 349400
rect 475200 347400 478600 348000
rect 475200 346000 475800 347400
rect 477200 346000 478600 347400
rect 475200 345400 478600 346000
rect 475200 344000 475800 345400
rect 477200 344000 478600 345400
rect 475200 343400 478600 344000
rect 475200 342000 475800 343400
rect 477200 342000 478600 343400
rect 475200 341400 478600 342000
rect 475200 340000 475800 341400
rect 477200 340000 478600 341400
rect 475200 339400 478600 340000
rect 475200 338000 475800 339400
rect 477200 338000 478600 339400
rect 475200 337400 478600 338000
rect 475200 336000 475800 337400
rect 477200 336000 478600 337400
rect 475200 335400 478600 336000
rect 475200 334000 475800 335400
rect 477200 334000 478600 335400
rect 475200 333400 478600 334000
rect 475200 332000 475800 333400
rect 477200 332000 478600 333400
rect 475200 331400 478600 332000
rect 475200 330000 475800 331400
rect 477200 330000 478600 331400
rect 475200 329400 478600 330000
rect 475200 328000 475800 329400
rect 477200 328000 478600 329400
rect 475200 327400 478600 328000
rect 475200 326000 475800 327400
rect 477200 326000 478600 327400
rect 475200 325400 478600 326000
rect 475200 324000 475800 325400
rect 477200 324000 478600 325400
rect 475200 323400 478600 324000
rect 475200 322000 475800 323400
rect 477200 322000 478600 323400
rect 475200 321400 478600 322000
rect 475200 320000 475800 321400
rect 477200 320000 478600 321400
rect 475200 319400 478600 320000
rect 475200 318000 475800 319400
rect 477200 318000 478600 319400
rect 475200 317400 478600 318000
rect 475200 316000 475800 317400
rect 477200 316000 478600 317400
rect 475200 315400 478600 316000
rect 475200 314000 475800 315400
rect 477200 314000 478600 315400
rect 475200 313400 478600 314000
rect 475200 312000 475800 313400
rect 477200 312000 478600 313400
rect 475200 311400 478600 312000
rect 475200 310000 475800 311400
rect 477200 310000 478600 311400
rect 475200 309400 478600 310000
rect 475200 308000 475800 309400
rect 477200 308000 478600 309400
rect 475200 307400 478600 308000
rect 475200 306000 475800 307400
rect 477200 306000 478600 307400
rect 475200 305400 478600 306000
rect 475200 304000 475800 305400
rect 477200 304000 478600 305400
rect 475200 303400 478600 304000
rect 475200 302000 475800 303400
rect 477200 302000 478600 303400
rect 475200 301400 478600 302000
rect 475200 300000 475800 301400
rect 477200 300000 478600 301400
rect 475200 299400 478600 300000
rect 475200 298000 475800 299400
rect 477200 298000 478600 299400
rect 475200 297400 478600 298000
rect 475200 296000 475800 297400
rect 477200 296000 478600 297400
rect 475200 295400 478600 296000
rect 475200 294000 475800 295400
rect 477200 294000 478600 295400
rect 475200 293400 478600 294000
rect 475200 292000 475800 293400
rect 477200 292000 478600 293400
rect 475200 291400 478600 292000
rect 475200 290000 475800 291400
rect 477200 290000 478600 291400
rect 475200 289400 478600 290000
rect 475200 288000 475800 289400
rect 477200 288000 478600 289400
rect 475200 287400 478600 288000
rect 475200 286000 475800 287400
rect 477200 286000 478600 287400
rect 475200 285400 478600 286000
rect 475200 284000 475800 285400
rect 477200 284000 478600 285400
rect 475200 283400 478600 284000
rect 475200 282000 475800 283400
rect 477200 282000 478600 283400
rect 475200 281400 478600 282000
rect 475200 280000 475800 281400
rect 477200 280000 478600 281400
rect 475200 279400 478600 280000
rect 475200 278000 475800 279400
rect 477200 278000 478600 279400
rect 475200 277400 478600 278000
rect 475200 276000 475800 277400
rect 477200 276000 478600 277400
rect 475200 275400 478600 276000
rect 475200 274000 475800 275400
rect 477200 274000 478600 275400
rect 475200 273400 478600 274000
rect 475200 272000 475800 273400
rect 477200 272000 478600 273400
rect 475200 271400 478600 272000
rect 475200 270000 475800 271400
rect 477200 270000 478600 271400
rect 475200 269400 478600 270000
rect 475200 268000 475800 269400
rect 477200 268000 478600 269400
rect 475200 267400 478600 268000
rect 475200 266000 475800 267400
rect 477200 266000 478600 267400
rect 475200 265400 478600 266000
rect 475200 264000 475800 265400
rect 477200 264000 478600 265400
rect 475200 263400 478600 264000
rect 475200 262000 475800 263400
rect 477200 262000 478600 263400
rect 475200 261400 478600 262000
rect 475200 260000 475800 261400
rect 477200 260000 478600 261400
rect 475200 259400 478600 260000
rect 475200 258000 475800 259400
rect 477200 258000 478600 259400
rect 475200 257400 478600 258000
rect 475200 256000 475800 257400
rect 477200 256000 478600 257400
rect 475200 255400 478600 256000
rect 475200 254000 475800 255400
rect 477200 254000 478600 255400
rect 475200 253400 478600 254000
rect 475200 252000 475800 253400
rect 477200 252000 478600 253400
rect 475200 251400 478600 252000
rect 475200 250000 475800 251400
rect 477200 250000 478600 251400
rect 475200 249400 478600 250000
rect 475200 248000 475800 249400
rect 477200 248000 478600 249400
rect 475200 247400 478600 248000
rect 475200 246000 475800 247400
rect 477200 246000 478600 247400
rect 475200 245400 478600 246000
rect 475200 244000 475800 245400
rect 477200 244000 478600 245400
rect 475200 243400 478600 244000
rect 475200 242000 475800 243400
rect 477200 242000 478600 243400
rect 475200 241400 478600 242000
rect 475200 240000 475800 241400
rect 477200 240000 478600 241400
rect 568600 241530 577600 242800
rect 568600 240370 568700 241530
rect 569770 241520 577600 241530
rect 577420 240400 577600 241520
rect 576370 240370 577600 240400
rect 568600 240000 577600 240370
rect 475200 239400 478600 240000
rect 475200 238000 475800 239400
rect 477200 238000 478600 239400
rect 475200 237400 478600 238000
rect 475200 236000 475800 237400
rect 477200 236000 478600 237400
rect 475200 235400 478600 236000
rect 475200 234000 475800 235400
rect 477200 234000 478600 235400
rect 475200 233400 478600 234000
rect 475200 232000 475800 233400
rect 477200 232000 478600 233400
rect 475200 231400 478600 232000
rect 475200 230000 475800 231400
rect 477200 230000 478600 231400
rect 475200 229400 478600 230000
rect 475200 228000 475800 229400
rect 477200 228000 478600 229400
rect 475200 227400 478600 228000
rect 475200 226000 475800 227400
rect 477200 226000 478600 227400
rect 475200 225400 478600 226000
rect 475200 224000 475800 225400
rect 477200 224000 478600 225400
rect 475200 223400 478600 224000
rect 475200 222000 475800 223400
rect 477200 222000 478600 223400
rect 475200 221400 478600 222000
rect 475200 220000 475800 221400
rect 477200 220000 478600 221400
rect 475200 219400 478600 220000
rect 475200 218000 475800 219400
rect 477200 218000 478600 219400
rect 475200 217400 478600 218000
rect 475200 216000 475800 217400
rect 477200 216000 478600 217400
rect 475200 215400 478600 216000
rect 475200 214000 475800 215400
rect 477200 214000 478600 215400
rect 475200 213400 478600 214000
rect 475200 212000 475800 213400
rect 477200 212000 478600 213400
rect 475200 211400 478600 212000
rect 475200 210000 475800 211400
rect 477200 210000 478600 211400
rect 475200 209400 478600 210000
rect 475200 208000 475800 209400
rect 477200 208000 478600 209400
rect 475200 207400 478600 208000
rect 475200 206000 475800 207400
rect 477200 206000 478600 207400
rect 475200 205400 478600 206000
rect 475200 204000 475800 205400
rect 477200 204000 478600 205400
rect 475200 203400 478600 204000
rect 475200 202000 475800 203400
rect 477200 202000 478600 203400
rect 475200 201400 478600 202000
rect 475200 200000 475800 201400
rect 477200 200000 478600 201400
rect 475200 199400 478600 200000
rect 475200 198000 475800 199400
rect 477200 198000 478600 199400
rect 475200 197400 478600 198000
rect 475200 196000 475800 197400
rect 477200 196000 478600 197400
rect 475200 195400 478600 196000
rect 475200 194000 475800 195400
rect 477200 194000 478600 195400
rect 475200 193400 478600 194000
rect 475200 192000 475800 193400
rect 477200 192000 478600 193400
rect 475200 191400 478600 192000
rect 475200 190000 475800 191400
rect 477200 190000 478600 191400
rect 475200 189400 478600 190000
rect 579200 201000 581200 201200
rect 579200 198160 579460 201000
rect 580960 198160 581200 201000
rect 579200 189900 579500 198160
rect 580900 189900 581200 198160
rect 579200 189500 581200 189900
rect 475200 188000 475800 189400
rect 477200 188000 478600 189400
rect 475200 187400 478600 188000
rect 475200 186000 475800 187400
rect 477200 186000 478600 187400
rect 475200 185400 478600 186000
rect 475200 184000 475800 185400
rect 477200 184000 478600 185400
rect 475200 183400 478600 184000
rect 475200 182000 475800 183400
rect 477200 182000 478600 183400
rect 475200 181400 478600 182000
rect 475200 180000 475800 181400
rect 477200 180000 478600 181400
rect 475200 179400 478600 180000
rect 475200 178000 475800 179400
rect 477200 178000 478600 179400
rect 475200 177400 478600 178000
rect 475200 176000 475800 177400
rect 477200 176000 478600 177400
rect 475200 175400 478600 176000
rect 576260 175800 579530 175830
rect 475200 174000 475800 175400
rect 477200 174000 478600 175400
rect 475200 173400 478600 174000
rect 475200 172000 475800 173400
rect 477200 172000 478600 173400
rect 475200 171400 478600 172000
rect 475200 170000 475800 171400
rect 477200 170000 478600 171400
rect 475200 169400 478600 170000
rect 475200 168000 475800 169400
rect 477200 168000 478600 169400
rect 475200 167400 478600 168000
rect 475200 166000 475800 167400
rect 477200 166000 478600 167400
rect 576200 175500 579600 175800
rect 576200 167200 576400 175500
rect 579400 167200 579600 175500
rect 576200 166600 579600 167200
rect 475200 165400 478600 166000
rect 475200 164000 475800 165400
rect 477200 164000 478600 165400
rect 475200 163400 478600 164000
rect 475200 162000 475800 163400
rect 477200 162000 478600 163400
rect 475200 161400 478600 162000
rect 475200 160000 475800 161400
rect 477200 160000 478600 161400
rect 475200 159400 478600 160000
rect 475200 158000 475800 159400
rect 477200 158000 478600 159400
rect 475200 157400 478600 158000
rect 475200 156000 475800 157400
rect 477200 156000 478600 157400
rect 475200 155400 478600 156000
rect 475200 154000 475800 155400
rect 477200 154000 478600 155400
rect 475200 153400 478600 154000
rect 475200 152000 475800 153400
rect 477200 152000 478600 153400
rect 572960 152600 576640 152630
rect 475200 151400 478600 152000
rect 475200 150000 475800 151400
rect 477200 150000 478600 151400
rect 475200 149400 478600 150000
rect 475200 148000 475800 149400
rect 477200 148000 478600 149400
rect 475200 147400 478600 148000
rect 475200 146000 475800 147400
rect 477200 146000 478600 147400
rect 475200 145400 478600 146000
rect 475200 144000 475800 145400
rect 477200 144000 478600 145400
rect 475200 143400 478600 144000
rect 475200 142000 475800 143400
rect 477200 142000 478600 143400
rect 572900 152000 576700 152600
rect 572900 151830 573200 152000
rect 572900 148990 573150 151830
rect 572900 143700 573200 148990
rect 576200 143700 576700 152000
rect 572900 143300 576700 143700
rect 475200 141400 478600 142000
rect 475200 140000 475800 141400
rect 477200 140000 478600 141400
rect 475200 139400 478600 140000
rect 475200 138000 475800 139400
rect 477200 138000 478600 139400
rect 475200 137400 478600 138000
rect 475200 136000 475800 137400
rect 477200 136000 478600 137400
rect 475200 135400 478600 136000
rect 475200 134000 475800 135400
rect 477200 134000 478600 135400
rect 475200 133400 478600 134000
rect 475200 132000 475800 133400
rect 477200 132000 478600 133400
rect 475200 131400 478600 132000
rect 475200 130000 475800 131400
rect 477200 130000 478600 131400
rect 475200 129400 478600 130000
rect 475200 128000 475800 129400
rect 477200 128000 478600 129400
rect 475200 127400 478600 128000
rect 475200 126000 475800 127400
rect 477200 126000 478600 127400
rect 475200 125400 478600 126000
rect 475200 124000 475800 125400
rect 477200 124000 478600 125400
rect 475200 123400 478600 124000
rect 475200 122000 475800 123400
rect 477200 122000 478600 123400
rect 570290 130770 578040 131480
rect 570290 123400 570850 130770
rect 577320 123400 578040 130770
rect 570290 123020 578040 123400
rect 475200 121400 478600 122000
rect 475200 120000 475800 121400
rect 477200 120000 478600 121400
rect 475200 119400 478600 120000
rect 475200 118000 475800 119400
rect 477200 118000 478600 119400
rect 475200 117400 478600 118000
rect 475200 116000 475800 117400
rect 477200 116000 478600 117400
rect 475200 115400 478600 116000
rect 475200 114000 475800 115400
rect 477200 114000 478600 115400
rect 475200 113400 478600 114000
rect 475200 112000 475800 113400
rect 477200 112000 478600 113400
rect 475200 111400 478600 112000
rect 475200 110000 475800 111400
rect 477200 110000 478600 111400
rect 475200 109400 478600 110000
rect 475200 108000 475800 109400
rect 477200 108000 478600 109400
rect 475200 107400 478600 108000
rect 475200 106000 475800 107400
rect 477200 106000 478600 107400
rect 475200 105400 478600 106000
rect 475200 104000 475800 105400
rect 477200 104000 478600 105400
rect 475200 103400 478600 104000
rect 475200 102000 475800 103400
rect 477200 102000 478600 103400
rect 475200 101400 478600 102000
rect 475200 100000 475800 101400
rect 477200 100000 478600 101400
rect 475200 99400 478600 100000
rect 475200 98000 475800 99400
rect 477200 98000 478600 99400
rect 475200 97400 478600 98000
rect 475200 96000 475800 97400
rect 477200 96000 478600 97400
rect 475200 95400 478600 96000
rect 475200 94000 475800 95400
rect 477200 94000 478600 95400
rect 475200 93400 478600 94000
rect 475200 92000 475800 93400
rect 477200 92000 478600 93400
rect 475200 91400 478600 92000
rect 475200 90000 475800 91400
rect 477200 90000 478600 91400
rect 475200 89400 478600 90000
rect 475200 88000 475800 89400
rect 477200 88000 478600 89400
rect 475200 87400 478600 88000
rect 475200 86000 475800 87400
rect 477200 86000 478600 87400
rect 475200 85400 478600 86000
rect 475200 84000 475800 85400
rect 477200 84000 478600 85400
rect 475200 83400 478600 84000
rect 475200 82000 475800 83400
rect 477200 82000 478600 83400
rect 475200 81400 478600 82000
rect 475200 80000 475800 81400
rect 477200 80000 478600 81400
rect 475200 79400 478600 80000
rect 475200 78000 475800 79400
rect 477200 78000 478600 79400
rect 475200 77400 478600 78000
rect 475200 76000 475800 77400
rect 477200 76000 478600 77400
rect 475200 75400 478600 76000
rect 475200 74000 475800 75400
rect 477200 74000 478600 75400
rect 475200 73400 478600 74000
rect 475200 72000 475800 73400
rect 477200 72000 478600 73400
rect 475200 71400 478600 72000
rect 475200 70000 475800 71400
rect 477200 70000 478600 71400
rect 475200 69400 478600 70000
rect 475200 68000 475800 69400
rect 477200 68000 478600 69400
rect 475200 67400 478600 68000
rect 475200 66000 475800 67400
rect 477200 66000 478600 67400
rect 475200 65400 478600 66000
rect 475200 64000 475800 65400
rect 477200 64000 478600 65400
rect 475200 63400 478600 64000
rect 475200 62000 475800 63400
rect 477200 62000 478600 63400
rect 475200 61400 478600 62000
rect 475200 60000 475800 61400
rect 477200 60000 478600 61400
rect 475200 59400 478600 60000
rect 475200 58000 475800 59400
rect 477200 58000 478600 59400
rect 475200 57400 478600 58000
rect 475200 56000 475800 57400
rect 477200 56000 478600 57400
rect 475200 55400 478600 56000
rect 475200 54000 475800 55400
rect 477200 54000 478600 55400
rect 475200 53400 478600 54000
rect 475200 52000 475800 53400
rect 477200 52000 478600 53400
rect 475200 51400 478600 52000
rect 475200 50000 475800 51400
rect 477200 50000 478600 51400
rect 475200 49400 478600 50000
rect 475200 48000 475800 49400
rect 477200 48000 478600 49400
rect 475200 47400 478600 48000
rect 475200 46000 475800 47400
rect 477200 46000 478600 47400
rect 475200 45400 478600 46000
rect 475200 44000 475800 45400
rect 477200 44000 478600 45400
rect 475200 43400 478600 44000
rect 475200 42000 475800 43400
rect 477200 42000 478600 43400
rect 475200 41400 478600 42000
rect 475200 40000 475800 41400
rect 477200 40000 478600 41400
rect 475200 39400 478600 40000
rect 475200 38000 475800 39400
rect 477200 38000 478600 39400
rect 475200 37400 478600 38000
rect 475200 36000 475800 37400
rect 477200 36000 478600 37400
rect 475200 35400 478600 36000
rect 475200 34000 475800 35400
rect 477200 34000 478600 35400
rect 475200 33400 478600 34000
rect 475200 32000 475800 33400
rect 477200 32000 478600 33400
rect 475200 31400 478600 32000
rect 475200 30000 475800 31400
rect 477200 30000 478600 31400
rect 475200 29400 478600 30000
rect 475200 28000 475800 29400
rect 477200 28000 478600 29400
rect 475200 27400 478600 28000
rect 475200 26000 475800 27400
rect 477200 26000 478600 27400
rect 475200 25400 478600 26000
rect 475200 24000 475800 25400
rect 477200 24000 478600 25400
rect 475200 23400 478600 24000
rect 475200 22000 475800 23400
rect 477200 22000 478600 23400
rect 475200 21400 478600 22000
rect 475200 20000 475800 21400
rect 477200 20000 478600 21400
rect 475200 19400 478600 20000
rect 475200 18000 475800 19400
rect 477200 18000 478600 19400
rect 475200 17400 478600 18000
rect 475200 16000 475800 17400
rect 477200 16000 478600 17400
rect 475200 15400 478600 16000
rect 475200 14000 475800 15400
rect 477200 14000 478600 15400
rect 475200 13400 478600 14000
rect 475200 12000 475800 13400
rect 477200 12000 478600 13400
rect 475200 11400 478600 12000
rect 475200 10000 475800 11400
rect 477200 10000 478600 11400
rect 475200 9400 478600 10000
rect 475200 8000 475800 9400
rect 477200 8000 478600 9400
rect 475200 7400 478600 8000
rect 475200 6000 475800 7400
rect 477200 6000 478600 7400
rect 475200 5400 478600 6000
rect 475200 4400 475800 5400
rect 15800 4000 475800 4400
rect 477200 4400 478600 5400
rect 477200 4000 568600 4400
rect 15800 2200 568600 4000
rect 475200 2000 478600 2200
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sky130_ef_io__bare_pad  BarePad_0
timestamp 1661870102
transform 1 0 569940 0 1 242260
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_1
timestamp 1661870102
transform 1 0 570860 0 1 187820
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_2
timestamp 1661870102
transform 1 0 570860 0 1 164820
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_3
timestamp 1661870102
transform 1 0 570860 0 1 141820
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_4
timestamp 1661870102
transform 1 0 570860 0 1 118820
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_5
timestamp 1661870102
transform 0 -1 528670 1 0 493270
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_6
timestamp 1661870102
transform 0 -1 528670 1 0 470270
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_7
timestamp 1661870102
transform 0 -1 551670 1 0 470270
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_8
timestamp 1661870102
transform 0 -1 574670 1 0 470270
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_9
timestamp 1661870102
transform -1 0 551420 0 -1 532090
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_10
timestamp 1661870102
transform -1 0 574420 0 -1 532090
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_11
timestamp 1661870102
transform -1 0 574420 0 -1 555090
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_12
timestamp 1661870102
transform -1 0 574420 0 -1 578090
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_13
timestamp 1661870102
transform -1 0 498830 0 -1 531960
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_14
timestamp 1661870102
transform -1 0 521830 0 -1 531960
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_15
timestamp 1661870102
transform -1 0 521830 0 -1 554960
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_16
timestamp 1661870102
transform -1 0 521830 0 -1 577960
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_17
timestamp 1661870102
transform -1 0 506820 0 -1 627620
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_18
timestamp 1661870102
transform -1 0 529820 0 -1 627620
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_19
timestamp 1661870102
transform -1 0 529820 0 -1 650620
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  BarePad_20
timestamp 1661870102
transform -1 0 529820 0 -1 673620
box -540 -540 12540 14540
use ComparatorQpixLayout  ComparatorQpixLayout_0
timestamp 1663612738
transform 0 -1 6052 1 0 525380
box 1330 -4580 8130 180
use RingOsl_v0_3stage  RingOsl_v0_3stage_1
timestamp 1663601856
transform 0 -1 577480 1 0 354470
box -740 -720 7730 2330
use classic-opamp  classic-opamp_0
timestamp 1663455834
transform 0 -1 573160 1 0 209510
box -5040 -7950 5960 250
use classic-opamp  classic-opamp_1
timestamp 1663455834
transform -1 0 561420 0 -1 496490
box -5040 -7950 5960 250
use classic-opamp  classic-opamp_2
timestamp 1663455834
transform 0 1 548200 -1 0 564840
box -5040 -7950 5960 250
use classic-opamp  classic-opamp_3
timestamp 1663455834
transform 0 1 495610 -1 0 564710
box -5040 -7950 5960 250
use classic-opamp  classic-opamp_4
timestamp 1663455834
transform 0 1 503600 -1 0 660370
box -5040 -7950 5960 250
use classic-opamp  classic-opamp_5
timestamp 1663455834
transform 0 -1 6193 1 0 336580
box -5040 -7950 5960 250
use mosarray  mosarray_0
timestamp 1663665281
transform 1 0 3180 0 1 3240
box 13000 -250 564910 675000
use opamp_diego  opamp_diego_0
timestamp 1606921152
transform 0 -1 571589 1 0 213341
box 2069 -10028 26971 3199
use opamp_diego  opamp_diego_1
timestamp 1606921152
transform -1 0 557589 0 -1 495969
box 2069 -10028 26971 3199
use opamp_diego  opamp_diego_2
timestamp 1606921152
transform 0 1 548721 -1 0 561009
box 2069 -10028 26971 3199
use opamp_diego  opamp_diego_3
timestamp 1606921152
transform 0 1 496131 -1 0 560879
box 2069 -10028 26971 3199
use opamp_diego  opamp_diego_4
timestamp 1606921152
transform 0 1 504121 -1 0 656539
box 2069 -10028 26971 3199
use opamp_diego  opamp_diego_5
timestamp 1606921152
transform 0 -1 5672 1 0 340411
box 2069 -10028 26971 3199
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_0
timestamp 1662310366
transform 0 1 574941 -1 0 365251
box -38 -49 2150 715
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_1
timestamp 1662310366
transform 0 1 577741 -1 0 365251
box -38 -49 2150 715
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_2
timestamp 1662310366
transform 0 -1 8149 1 0 534649
box -38 -49 2150 715
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
