magic
tech sky130A
timestamp 1663655995
<< nwell >>
rect 55383 219286 57006 220939
rect 77883 219286 79506 220939
rect 100383 219286 102006 220939
rect 122883 219286 124506 220939
rect 145383 219286 147006 220939
rect 55383 196286 57006 197368
rect 77883 196286 79506 197368
rect 100383 196286 102006 197368
rect 122883 196286 124506 197368
rect 145383 196286 147006 197368
rect 55383 173286 57006 174368
rect 77883 173286 79506 174368
rect 100383 173286 102006 174368
rect 122883 173286 124506 174368
rect 145383 173286 147006 174368
rect 55383 150286 57006 151368
rect 77883 150286 79506 151368
rect 100383 150286 102006 151368
rect 122883 150286 124506 151368
rect 145383 150286 147006 151368
rect 55383 127286 57006 128368
rect 77883 127286 79506 128368
rect 100383 127286 102006 128368
rect 122883 127286 124506 128368
rect 145383 127286 147006 128368
rect 55383 104286 57006 105368
rect 77883 104286 79506 105368
rect 100383 104286 102006 105368
rect 122883 104286 124506 105368
rect 145383 104286 147006 105368
rect 55383 81286 57006 82368
rect 77883 81286 79506 82368
rect 100383 81286 102006 82368
rect 122883 81286 124506 82368
rect 145383 81286 147006 82368
rect 55383 58286 57006 59368
rect 77883 58286 79506 59368
rect 100383 58286 102006 59368
rect 122883 58286 124506 59368
rect 145383 58286 147006 59368
rect 55383 35286 57006 36368
rect 77883 35286 79506 36368
rect 100383 35286 102006 36368
rect 122883 35286 124506 36368
rect 145383 35286 147006 36368
rect 54912 2236 57618 13659
rect 77519 2236 80225 13659
rect 99885 2116 102591 13539
rect 122552 2236 125258 13659
rect 144979 2357 147685 13780
<< pmoslvt >>
rect 56156 220074 56191 220116
rect 78666 220074 78716 220116
rect 101166 220074 101266 220116
rect 123666 220074 123866 220116
rect 146166 220074 146566 220116
rect 56156 197061 56191 197116
rect 78666 197061 78716 197116
rect 101166 197061 101266 197116
rect 123666 197061 123866 197116
rect 146166 197061 146566 197116
rect 56156 174052 56191 174116
rect 78666 174052 78716 174116
rect 101166 174052 101266 174116
rect 123666 174052 123866 174116
rect 146166 174052 146566 174116
rect 56156 151032 56191 151116
rect 78666 151032 78716 151116
rect 101166 151032 101266 151116
rect 123666 151032 123866 151116
rect 146166 151032 146566 151116
rect 56156 128016 56191 128116
rect 78666 128016 78716 128116
rect 101166 128016 101266 128116
rect 123666 128016 123866 128116
rect 146166 128016 146566 128116
rect 56156 104951 56191 105116
rect 78666 104951 78716 105116
rect 101166 104951 101266 105116
rect 123666 104951 123866 105116
rect 146166 104951 146566 105116
rect 56156 81816 56191 82116
rect 78666 81816 78716 82116
rect 101166 81816 101266 82116
rect 123666 81816 123866 82116
rect 146166 81816 146566 82116
rect 56156 58616 56191 59116
rect 78666 58616 78716 59116
rect 101166 58616 101266 59116
rect 123666 58616 123866 59116
rect 146166 58616 146566 59116
rect 56156 35416 56191 36116
rect 78666 35416 78716 36116
rect 101166 35416 101266 36116
rect 123666 35416 123866 36116
rect 146166 35416 146566 36116
rect 56156 3116 56191 13116
rect 78666 3116 78716 13116
rect 101166 3116 101266 13116
rect 123666 3116 123866 13116
rect 146166 3116 146566 13116
<< pdiff >>
rect 56056 220103 56156 220116
rect 56056 220086 56068 220103
rect 56144 220086 56156 220103
rect 56056 220074 56156 220086
rect 56191 220103 56291 220116
rect 56191 220086 56203 220103
rect 56279 220086 56291 220103
rect 56191 220074 56291 220086
rect 78566 220103 78666 220116
rect 78566 220086 78578 220103
rect 78654 220086 78666 220103
rect 78566 220074 78666 220086
rect 78716 220103 78816 220116
rect 78716 220086 78728 220103
rect 78804 220086 78816 220103
rect 78716 220074 78816 220086
rect 101066 220103 101166 220116
rect 101066 220086 101078 220103
rect 101154 220086 101166 220103
rect 101066 220074 101166 220086
rect 101266 220103 101366 220116
rect 101266 220086 101278 220103
rect 101354 220086 101366 220103
rect 101266 220074 101366 220086
rect 123566 220103 123666 220116
rect 123566 220086 123578 220103
rect 123654 220086 123666 220103
rect 123566 220074 123666 220086
rect 123866 220103 123966 220116
rect 123866 220086 123878 220103
rect 123954 220086 123966 220103
rect 123866 220074 123966 220086
rect 146066 220103 146166 220116
rect 146066 220086 146078 220103
rect 146154 220086 146166 220103
rect 146066 220074 146166 220086
rect 146566 220103 146666 220116
rect 146566 220086 146578 220103
rect 146654 220086 146666 220103
rect 146566 220074 146666 220086
rect 56056 197103 56156 197116
rect 56056 197073 56068 197103
rect 56144 197073 56156 197103
rect 56056 197061 56156 197073
rect 56191 197103 56291 197116
rect 56191 197073 56203 197103
rect 56279 197073 56291 197103
rect 56191 197061 56291 197073
rect 78566 197103 78666 197116
rect 78566 197073 78578 197103
rect 78654 197073 78666 197103
rect 78566 197061 78666 197073
rect 78716 197103 78816 197116
rect 78716 197073 78728 197103
rect 78804 197073 78816 197103
rect 78716 197061 78816 197073
rect 101066 197103 101166 197116
rect 101066 197073 101078 197103
rect 101154 197073 101166 197103
rect 101066 197061 101166 197073
rect 101266 197103 101366 197116
rect 101266 197073 101278 197103
rect 101354 197073 101366 197103
rect 101266 197061 101366 197073
rect 123566 197103 123666 197116
rect 123566 197073 123578 197103
rect 123654 197073 123666 197103
rect 123566 197061 123666 197073
rect 123866 197103 123966 197116
rect 123866 197073 123878 197103
rect 123954 197073 123966 197103
rect 123866 197061 123966 197073
rect 146066 197103 146166 197116
rect 146066 197073 146078 197103
rect 146154 197073 146166 197103
rect 146066 197061 146166 197073
rect 146566 197103 146666 197116
rect 146566 197073 146578 197103
rect 146654 197073 146666 197103
rect 146566 197061 146666 197073
rect 56056 174103 56156 174116
rect 56056 174064 56068 174103
rect 56144 174064 56156 174103
rect 56056 174052 56156 174064
rect 56191 174103 56291 174116
rect 56191 174064 56203 174103
rect 56279 174064 56291 174103
rect 56191 174052 56291 174064
rect 78566 174103 78666 174116
rect 78566 174064 78578 174103
rect 78654 174064 78666 174103
rect 78566 174052 78666 174064
rect 78716 174103 78816 174116
rect 78716 174064 78728 174103
rect 78804 174064 78816 174103
rect 78716 174052 78816 174064
rect 101066 174103 101166 174116
rect 101066 174064 101078 174103
rect 101154 174064 101166 174103
rect 101066 174052 101166 174064
rect 101266 174103 101366 174116
rect 101266 174064 101278 174103
rect 101354 174064 101366 174103
rect 101266 174052 101366 174064
rect 123566 174103 123666 174116
rect 123566 174064 123578 174103
rect 123654 174064 123666 174103
rect 123566 174052 123666 174064
rect 123866 174103 123966 174116
rect 123866 174064 123878 174103
rect 123954 174064 123966 174103
rect 123866 174052 123966 174064
rect 146066 174103 146166 174116
rect 146066 174064 146078 174103
rect 146154 174064 146166 174103
rect 146066 174052 146166 174064
rect 146566 174103 146666 174116
rect 146566 174064 146578 174103
rect 146654 174064 146666 174103
rect 146566 174052 146666 174064
rect 56056 151103 56156 151116
rect 56056 151044 56068 151103
rect 56144 151044 56156 151103
rect 56056 151032 56156 151044
rect 56191 151103 56291 151116
rect 56191 151044 56203 151103
rect 56279 151044 56291 151103
rect 56191 151032 56291 151044
rect 78566 151103 78666 151116
rect 78566 151044 78578 151103
rect 78654 151044 78666 151103
rect 78566 151032 78666 151044
rect 78716 151103 78816 151116
rect 78716 151044 78728 151103
rect 78804 151044 78816 151103
rect 78716 151032 78816 151044
rect 101066 151103 101166 151116
rect 101066 151044 101078 151103
rect 101154 151044 101166 151103
rect 101066 151032 101166 151044
rect 101266 151103 101366 151116
rect 101266 151044 101278 151103
rect 101354 151044 101366 151103
rect 101266 151032 101366 151044
rect 123566 151103 123666 151116
rect 123566 151044 123578 151103
rect 123654 151044 123666 151103
rect 123566 151032 123666 151044
rect 123866 151103 123966 151116
rect 123866 151044 123878 151103
rect 123954 151044 123966 151103
rect 123866 151032 123966 151044
rect 146066 151103 146166 151116
rect 146066 151044 146078 151103
rect 146154 151044 146166 151103
rect 146066 151032 146166 151044
rect 146566 151103 146666 151116
rect 146566 151044 146578 151103
rect 146654 151044 146666 151103
rect 146566 151032 146666 151044
rect 56056 128103 56156 128116
rect 56056 128028 56068 128103
rect 56144 128028 56156 128103
rect 56056 128016 56156 128028
rect 56191 128103 56291 128116
rect 56191 128028 56203 128103
rect 56279 128028 56291 128103
rect 56191 128016 56291 128028
rect 78566 128103 78666 128116
rect 78566 128028 78578 128103
rect 78654 128028 78666 128103
rect 78566 128016 78666 128028
rect 78716 128103 78816 128116
rect 78716 128028 78728 128103
rect 78804 128028 78816 128103
rect 78716 128016 78816 128028
rect 101066 128103 101166 128116
rect 101066 128028 101078 128103
rect 101154 128028 101166 128103
rect 101066 128016 101166 128028
rect 101266 128103 101366 128116
rect 101266 128028 101278 128103
rect 101354 128028 101366 128103
rect 101266 128016 101366 128028
rect 123566 128103 123666 128116
rect 123566 128028 123578 128103
rect 123654 128028 123666 128103
rect 123566 128016 123666 128028
rect 123866 128103 123966 128116
rect 123866 128028 123878 128103
rect 123954 128028 123966 128103
rect 123866 128016 123966 128028
rect 146066 128103 146166 128116
rect 146066 128028 146078 128103
rect 146154 128028 146166 128103
rect 146066 128016 146166 128028
rect 146566 128103 146666 128116
rect 146566 128028 146578 128103
rect 146654 128028 146666 128103
rect 146566 128016 146666 128028
rect 56056 105103 56156 105116
rect 56056 104963 56068 105103
rect 56144 104963 56156 105103
rect 56056 104951 56156 104963
rect 56191 105103 56291 105116
rect 56191 104963 56203 105103
rect 56279 104963 56291 105103
rect 56191 104951 56291 104963
rect 78566 105103 78666 105116
rect 78566 104963 78578 105103
rect 78654 104963 78666 105103
rect 78566 104951 78666 104963
rect 78716 105103 78816 105116
rect 78716 104963 78728 105103
rect 78804 104963 78816 105103
rect 78716 104951 78816 104963
rect 101066 105103 101166 105116
rect 101066 104963 101078 105103
rect 101154 104963 101166 105103
rect 101066 104951 101166 104963
rect 101266 105103 101366 105116
rect 101266 104963 101278 105103
rect 101354 104963 101366 105103
rect 101266 104951 101366 104963
rect 123566 105103 123666 105116
rect 123566 104963 123578 105103
rect 123654 104963 123666 105103
rect 123566 104951 123666 104963
rect 123866 105103 123966 105116
rect 123866 104963 123878 105103
rect 123954 104963 123966 105103
rect 123866 104951 123966 104963
rect 146066 105103 146166 105116
rect 146066 104963 146078 105103
rect 146154 104963 146166 105103
rect 146066 104951 146166 104963
rect 146566 105103 146666 105116
rect 146566 104963 146578 105103
rect 146654 104963 146666 105103
rect 146566 104951 146666 104963
rect 56056 82103 56156 82116
rect 56056 81828 56068 82103
rect 56144 81828 56156 82103
rect 56056 81816 56156 81828
rect 56191 82103 56291 82116
rect 56191 81828 56203 82103
rect 56279 81828 56291 82103
rect 56191 81816 56291 81828
rect 78566 82103 78666 82116
rect 78566 81828 78578 82103
rect 78654 81828 78666 82103
rect 78566 81816 78666 81828
rect 78716 82103 78816 82116
rect 78716 81828 78728 82103
rect 78804 81828 78816 82103
rect 78716 81816 78816 81828
rect 101066 82103 101166 82116
rect 101066 81828 101078 82103
rect 101154 81828 101166 82103
rect 101066 81816 101166 81828
rect 101266 82103 101366 82116
rect 101266 81828 101278 82103
rect 101354 81828 101366 82103
rect 101266 81816 101366 81828
rect 123566 82103 123666 82116
rect 123566 81828 123578 82103
rect 123654 81828 123666 82103
rect 123566 81816 123666 81828
rect 123866 82103 123966 82116
rect 123866 81828 123878 82103
rect 123954 81828 123966 82103
rect 123866 81816 123966 81828
rect 146066 82103 146166 82116
rect 146066 81828 146078 82103
rect 146154 81828 146166 82103
rect 146066 81816 146166 81828
rect 146566 82103 146666 82116
rect 146566 81828 146578 82103
rect 146654 81828 146666 82103
rect 146566 81816 146666 81828
rect 56056 59103 56156 59116
rect 56056 58628 56068 59103
rect 56144 58628 56156 59103
rect 56056 58616 56156 58628
rect 56191 59103 56291 59116
rect 56191 58628 56203 59103
rect 56279 58628 56291 59103
rect 56191 58616 56291 58628
rect 78566 59103 78666 59116
rect 78566 58628 78578 59103
rect 78654 58628 78666 59103
rect 78566 58616 78666 58628
rect 78716 59103 78816 59116
rect 78716 58628 78728 59103
rect 78804 58628 78816 59103
rect 78716 58616 78816 58628
rect 101066 59103 101166 59116
rect 101066 58628 101078 59103
rect 101154 58628 101166 59103
rect 101066 58616 101166 58628
rect 101266 59103 101366 59116
rect 101266 58628 101278 59103
rect 101354 58628 101366 59103
rect 101266 58616 101366 58628
rect 123566 59103 123666 59116
rect 123566 58628 123578 59103
rect 123654 58628 123666 59103
rect 123566 58616 123666 58628
rect 123866 59103 123966 59116
rect 123866 58628 123878 59103
rect 123954 58628 123966 59103
rect 146066 59103 146166 59116
rect 123866 58616 123966 58628
rect 146066 58628 146078 59103
rect 146154 58628 146166 59103
rect 146066 58616 146166 58628
rect 146566 59103 146666 59116
rect 146566 58628 146578 59103
rect 146654 58628 146666 59103
rect 146566 58616 146666 58628
rect 56056 36103 56156 36116
rect 56056 35428 56068 36103
rect 56144 35428 56156 36103
rect 56056 35416 56156 35428
rect 56191 36103 56291 36116
rect 56191 35428 56203 36103
rect 56279 35428 56291 36103
rect 56191 35416 56291 35428
rect 78566 36103 78666 36116
rect 78566 35428 78578 36103
rect 78654 35428 78666 36103
rect 78566 35416 78666 35428
rect 78716 36103 78816 36116
rect 78716 35428 78728 36103
rect 78804 35428 78816 36103
rect 78716 35416 78816 35428
rect 101066 36103 101166 36116
rect 101066 35428 101078 36103
rect 101154 35428 101166 36103
rect 101066 35416 101166 35428
rect 101266 36103 101366 36116
rect 101266 35428 101278 36103
rect 101354 35428 101366 36103
rect 101266 35416 101366 35428
rect 123566 36103 123666 36116
rect 123566 35428 123578 36103
rect 123654 35428 123666 36103
rect 123566 35416 123666 35428
rect 123866 36103 123966 36116
rect 123866 35428 123878 36103
rect 123954 35428 123966 36103
rect 123866 35416 123966 35428
rect 146066 36103 146166 36116
rect 146066 35428 146078 36103
rect 146154 35428 146166 36103
rect 146066 35416 146166 35428
rect 146566 36103 146666 36116
rect 146566 35428 146578 36103
rect 146654 35428 146666 36103
rect 146566 35416 146666 35428
rect 56056 13103 56156 13116
rect 56056 3128 56068 13103
rect 56144 3128 56156 13103
rect 56056 3116 56156 3128
rect 56191 13103 56291 13116
rect 56191 3128 56203 13103
rect 56279 3128 56291 13103
rect 56191 3116 56291 3128
rect 78566 13103 78666 13116
rect 78566 3128 78578 13103
rect 78654 3128 78666 13103
rect 78566 3116 78666 3128
rect 78716 13103 78816 13116
rect 78716 3128 78728 13103
rect 78804 3128 78816 13103
rect 78716 3116 78816 3128
rect 101066 13103 101166 13116
rect 101066 3128 101078 13103
rect 101154 3128 101166 13103
rect 101066 3116 101166 3128
rect 101266 13103 101366 13116
rect 101266 3128 101278 13103
rect 101354 3128 101366 13103
rect 101266 3116 101366 3128
rect 123566 13103 123666 13116
rect 123566 3128 123578 13103
rect 123654 3128 123666 13103
rect 123566 3116 123666 3128
rect 123866 13103 123966 13116
rect 123866 3128 123878 13103
rect 123954 3128 123966 13103
rect 123866 3116 123966 3128
rect 146066 13103 146166 13116
rect 146066 3128 146078 13103
rect 146154 3128 146166 13103
rect 146066 3116 146166 3128
rect 146566 13103 146666 13116
rect 146566 3128 146578 13103
rect 146654 3128 146666 13103
rect 146566 3116 146666 3128
<< pdiffc >>
rect 56068 220086 56144 220103
rect 56203 220086 56279 220103
rect 78578 220086 78654 220103
rect 78728 220086 78804 220103
rect 101078 220086 101154 220103
rect 101278 220086 101354 220103
rect 123578 220086 123654 220103
rect 123878 220086 123954 220103
rect 146078 220086 146154 220103
rect 146578 220086 146654 220103
rect 56068 197073 56144 197103
rect 56203 197073 56279 197103
rect 78578 197073 78654 197103
rect 78728 197073 78804 197103
rect 101078 197073 101154 197103
rect 101278 197073 101354 197103
rect 123578 197073 123654 197103
rect 123878 197073 123954 197103
rect 146078 197073 146154 197103
rect 146578 197073 146654 197103
rect 56068 174064 56144 174103
rect 56203 174064 56279 174103
rect 78578 174064 78654 174103
rect 78728 174064 78804 174103
rect 101078 174064 101154 174103
rect 101278 174064 101354 174103
rect 123578 174064 123654 174103
rect 123878 174064 123954 174103
rect 146078 174064 146154 174103
rect 146578 174064 146654 174103
rect 56068 151044 56144 151103
rect 56203 151044 56279 151103
rect 78578 151044 78654 151103
rect 78728 151044 78804 151103
rect 101078 151044 101154 151103
rect 101278 151044 101354 151103
rect 123578 151044 123654 151103
rect 123878 151044 123954 151103
rect 146078 151044 146154 151103
rect 146578 151044 146654 151103
rect 56068 128028 56144 128103
rect 56203 128028 56279 128103
rect 78578 128028 78654 128103
rect 78728 128028 78804 128103
rect 101078 128028 101154 128103
rect 101278 128028 101354 128103
rect 123578 128028 123654 128103
rect 123878 128028 123954 128103
rect 146078 128028 146154 128103
rect 146578 128028 146654 128103
rect 56068 104963 56144 105103
rect 56203 104963 56279 105103
rect 78578 104963 78654 105103
rect 78728 104963 78804 105103
rect 101078 104963 101154 105103
rect 101278 104963 101354 105103
rect 123578 104963 123654 105103
rect 123878 104963 123954 105103
rect 146078 104963 146154 105103
rect 146578 104963 146654 105103
rect 56068 81828 56144 82103
rect 56203 81828 56279 82103
rect 78578 81828 78654 82103
rect 78728 81828 78804 82103
rect 101078 81828 101154 82103
rect 101278 81828 101354 82103
rect 123578 81828 123654 82103
rect 123878 81828 123954 82103
rect 146078 81828 146154 82103
rect 146578 81828 146654 82103
rect 56068 58628 56144 59103
rect 56203 58628 56279 59103
rect 78578 58628 78654 59103
rect 78728 58628 78804 59103
rect 101078 58628 101154 59103
rect 101278 58628 101354 59103
rect 123578 58628 123654 59103
rect 123878 58628 123954 59103
rect 146078 58628 146154 59103
rect 146578 58628 146654 59103
rect 56068 35428 56144 36103
rect 56203 35428 56279 36103
rect 78578 35428 78654 36103
rect 78728 35428 78804 36103
rect 101078 35428 101154 36103
rect 101278 35428 101354 36103
rect 123578 35428 123654 36103
rect 123878 35428 123954 36103
rect 146078 35428 146154 36103
rect 146578 35428 146654 36103
rect 56068 3128 56144 13103
rect 56203 3128 56279 13103
rect 78578 3128 78654 13103
rect 78728 3128 78804 13103
rect 101078 3128 101154 13103
rect 101278 3128 101354 13103
rect 123578 3128 123654 13103
rect 123878 3128 123954 13103
rect 146078 3128 146154 13103
rect 146578 3128 146654 13103
<< nsubdiff >>
rect 55956 220103 56056 220116
rect 55956 220086 55969 220103
rect 56045 220086 56056 220103
rect 55956 220074 56056 220086
rect 78466 220103 78566 220116
rect 78466 220086 78479 220103
rect 78555 220086 78566 220103
rect 78466 220074 78566 220086
rect 100966 220103 101066 220116
rect 100966 220086 100979 220103
rect 101055 220086 101066 220103
rect 100966 220074 101066 220086
rect 123466 220103 123566 220116
rect 123466 220086 123479 220103
rect 123555 220086 123566 220103
rect 123466 220074 123566 220086
rect 145966 220103 146066 220116
rect 145966 220086 145979 220103
rect 146055 220086 146066 220103
rect 145966 220074 146066 220086
rect 55956 197103 56056 197116
rect 55956 197073 55969 197103
rect 56045 197073 56056 197103
rect 55956 197061 56056 197073
rect 78466 197103 78566 197116
rect 78466 197073 78479 197103
rect 78555 197073 78566 197103
rect 78466 197061 78566 197073
rect 100966 197103 101066 197116
rect 100966 197073 100979 197103
rect 101055 197073 101066 197103
rect 100966 197061 101066 197073
rect 123466 197103 123566 197116
rect 123466 197073 123479 197103
rect 123555 197073 123566 197103
rect 123466 197061 123566 197073
rect 145966 197103 146066 197116
rect 145966 197073 145979 197103
rect 146055 197073 146066 197103
rect 145966 197061 146066 197073
rect 55956 174103 56056 174116
rect 55956 174064 55969 174103
rect 56045 174064 56056 174103
rect 55956 174052 56056 174064
rect 78466 174103 78566 174116
rect 78466 174064 78479 174103
rect 78555 174064 78566 174103
rect 78466 174052 78566 174064
rect 100966 174103 101066 174116
rect 100966 174064 100979 174103
rect 101055 174064 101066 174103
rect 100966 174052 101066 174064
rect 123466 174103 123566 174116
rect 123466 174064 123479 174103
rect 123555 174064 123566 174103
rect 123466 174052 123566 174064
rect 145966 174103 146066 174116
rect 145966 174064 145979 174103
rect 146055 174064 146066 174103
rect 145966 174052 146066 174064
rect 55956 151103 56056 151116
rect 55956 151044 55969 151103
rect 56045 151044 56056 151103
rect 55956 151032 56056 151044
rect 78466 151103 78566 151116
rect 78466 151044 78479 151103
rect 78555 151044 78566 151103
rect 78466 151032 78566 151044
rect 100966 151103 101066 151116
rect 100966 151044 100979 151103
rect 101055 151044 101066 151103
rect 100966 151032 101066 151044
rect 123466 151103 123566 151116
rect 123466 151044 123479 151103
rect 123555 151044 123566 151103
rect 123466 151032 123566 151044
rect 145966 151103 146066 151116
rect 145966 151044 145979 151103
rect 146055 151044 146066 151103
rect 145966 151032 146066 151044
rect 55956 128103 56056 128116
rect 55956 128028 55969 128103
rect 56045 128028 56056 128103
rect 55956 128016 56056 128028
rect 78466 128103 78566 128116
rect 78466 128028 78479 128103
rect 78555 128028 78566 128103
rect 78466 128016 78566 128028
rect 100966 128103 101066 128116
rect 100966 128028 100979 128103
rect 101055 128028 101066 128103
rect 100966 128016 101066 128028
rect 123466 128103 123566 128116
rect 123466 128028 123479 128103
rect 123555 128028 123566 128103
rect 123466 128016 123566 128028
rect 145966 128103 146066 128116
rect 145966 128028 145979 128103
rect 146055 128028 146066 128103
rect 145966 128016 146066 128028
rect 55956 105103 56056 105116
rect 55956 104963 55969 105103
rect 56045 104963 56056 105103
rect 55956 104951 56056 104963
rect 78466 105103 78566 105116
rect 78466 104963 78479 105103
rect 78555 104963 78566 105103
rect 78466 104951 78566 104963
rect 100966 105103 101066 105116
rect 100966 104963 100979 105103
rect 101055 104963 101066 105103
rect 100966 104951 101066 104963
rect 123466 105103 123566 105116
rect 123466 104963 123479 105103
rect 123555 104963 123566 105103
rect 123466 104951 123566 104963
rect 145966 105103 146066 105116
rect 145966 104963 145979 105103
rect 146055 104963 146066 105103
rect 145966 104951 146066 104963
rect 55956 82103 56056 82116
rect 55956 81828 55969 82103
rect 56045 81828 56056 82103
rect 55956 81816 56056 81828
rect 78466 82103 78566 82116
rect 78466 81828 78479 82103
rect 78555 81828 78566 82103
rect 78466 81816 78566 81828
rect 100966 82103 101066 82116
rect 100966 81828 100979 82103
rect 101055 81828 101066 82103
rect 100966 81816 101066 81828
rect 123466 82103 123566 82116
rect 123466 81828 123479 82103
rect 123555 81828 123566 82103
rect 123466 81816 123566 81828
rect 145966 82103 146066 82116
rect 145966 81828 145979 82103
rect 146055 81828 146066 82103
rect 145966 81816 146066 81828
rect 55956 59103 56056 59116
rect 55956 58628 55969 59103
rect 56045 58628 56056 59103
rect 55956 58616 56056 58628
rect 78466 59103 78566 59116
rect 78466 58628 78479 59103
rect 78555 58628 78566 59103
rect 78466 58616 78566 58628
rect 100966 59103 101066 59116
rect 100966 58628 100979 59103
rect 101055 58628 101066 59103
rect 100966 58616 101066 58628
rect 123466 59103 123566 59116
rect 123466 58628 123479 59103
rect 123555 58628 123566 59103
rect 123466 58616 123566 58628
rect 145966 59103 146066 59116
rect 145966 58849 145979 59103
rect 145967 58628 145979 58849
rect 146055 58628 146066 59103
rect 145967 58616 146066 58628
rect 55956 36103 56056 36116
rect 55956 35428 55969 36103
rect 56045 35428 56056 36103
rect 55956 35416 56056 35428
rect 78466 36103 78566 36116
rect 78466 35428 78479 36103
rect 78555 35428 78566 36103
rect 78466 35416 78566 35428
rect 100966 36103 101066 36116
rect 100966 35428 100979 36103
rect 101055 35428 101066 36103
rect 100966 35416 101066 35428
rect 123466 36103 123566 36116
rect 123466 35428 123479 36103
rect 123555 35428 123566 36103
rect 123466 35416 123566 35428
rect 145966 36103 146066 36116
rect 145966 35428 145979 36103
rect 146055 35428 146066 36103
rect 145966 35416 146066 35428
rect 55956 13103 56056 13116
rect 55956 3128 55969 13103
rect 56045 3128 56056 13103
rect 55956 3116 56056 3128
rect 78466 13103 78566 13116
rect 78466 3128 78479 13103
rect 78555 3128 78566 13103
rect 78466 3116 78566 3128
rect 100966 13103 101066 13116
rect 100966 3128 100979 13103
rect 101055 3128 101066 13103
rect 100966 3116 101066 3128
rect 123466 13103 123566 13116
rect 123466 3128 123479 13103
rect 123555 3128 123566 13103
rect 123466 3116 123566 3128
rect 145966 13103 146066 13116
rect 145966 3128 145979 13103
rect 146055 3128 146066 13103
rect 145966 3116 146066 3128
<< nsubdiffcont >>
rect 55969 220086 56045 220103
rect 78479 220086 78555 220103
rect 100979 220086 101055 220103
rect 123479 220086 123555 220103
rect 145979 220086 146055 220103
rect 55969 197073 56045 197103
rect 78479 197073 78555 197103
rect 100979 197073 101055 197103
rect 123479 197073 123555 197103
rect 145979 197073 146055 197103
rect 55969 174064 56045 174103
rect 78479 174064 78555 174103
rect 100979 174064 101055 174103
rect 123479 174064 123555 174103
rect 145979 174064 146055 174103
rect 55969 151044 56045 151103
rect 78479 151044 78555 151103
rect 100979 151044 101055 151103
rect 123479 151044 123555 151103
rect 145979 151044 146055 151103
rect 55969 128028 56045 128103
rect 78479 128028 78555 128103
rect 100979 128028 101055 128103
rect 123479 128028 123555 128103
rect 145979 128028 146055 128103
rect 55969 104963 56045 105103
rect 78479 104963 78555 105103
rect 100979 104963 101055 105103
rect 123479 104963 123555 105103
rect 145979 104963 146055 105103
rect 55969 81828 56045 82103
rect 78479 81828 78555 82103
rect 100979 81828 101055 82103
rect 123479 81828 123555 82103
rect 145979 81828 146055 82103
rect 55969 58628 56045 59103
rect 78479 58628 78555 59103
rect 100979 58628 101055 59103
rect 123479 58628 123555 59103
rect 145979 58628 146055 59103
rect 55969 35428 56045 36103
rect 78479 35428 78555 36103
rect 100979 35428 101055 36103
rect 123479 35428 123555 36103
rect 145979 35428 146055 36103
rect 55969 3128 56045 13103
rect 78479 3128 78555 13103
rect 100979 3128 101055 13103
rect 123479 3128 123555 13103
rect 145979 3128 146055 13103
<< poly >>
rect 56139 220183 56199 220191
rect 56139 220149 56147 220183
rect 56191 220149 56199 220183
rect 56139 220141 56199 220149
rect 78649 220183 78716 220191
rect 78649 220149 78657 220183
rect 78691 220149 78716 220183
rect 78649 220141 78716 220149
rect 101149 220183 101199 220191
rect 101149 220149 101157 220183
rect 101191 220149 101199 220183
rect 101149 220141 101199 220149
rect 123649 220183 123866 220191
rect 123649 220149 123657 220183
rect 123860 220149 123866 220183
rect 123649 220141 123866 220149
rect 146149 220183 146566 220191
rect 146149 220149 146157 220183
rect 146149 220148 146178 220149
rect 146552 220148 146566 220183
rect 146149 220141 146566 220148
rect 56156 220116 56191 220141
rect 78666 220116 78716 220141
rect 101166 220116 101266 220141
rect 123666 220116 123866 220141
rect 146166 220116 146566 220141
rect 56156 220059 56191 220074
rect 78666 220059 78716 220074
rect 101166 220059 101266 220074
rect 123666 220059 123866 220074
rect 146166 220059 146566 220074
rect 56139 197183 56199 197191
rect 56139 197149 56147 197183
rect 56191 197149 56199 197183
rect 56139 197141 56199 197149
rect 78649 197183 78716 197191
rect 78649 197149 78657 197183
rect 78691 197149 78716 197183
rect 78649 197141 78716 197149
rect 101149 197183 101199 197191
rect 101149 197149 101157 197183
rect 101191 197149 101199 197183
rect 101149 197141 101199 197149
rect 123649 197183 123866 197191
rect 123649 197149 123657 197183
rect 123860 197149 123866 197183
rect 123649 197141 123866 197149
rect 146149 197183 146566 197191
rect 146149 197149 146157 197183
rect 146149 197148 146178 197149
rect 146552 197148 146566 197183
rect 146149 197141 146566 197148
rect 56156 197116 56191 197141
rect 78666 197116 78716 197141
rect 101166 197116 101266 197141
rect 123666 197116 123866 197141
rect 146166 197116 146566 197141
rect 56156 197048 56191 197061
rect 78666 197048 78716 197061
rect 101166 197047 101266 197061
rect 123666 197047 123866 197061
rect 146166 197047 146566 197061
rect 56139 174183 56199 174191
rect 56139 174149 56147 174183
rect 56191 174149 56199 174183
rect 56139 174141 56199 174149
rect 78649 174183 78716 174191
rect 78649 174149 78657 174183
rect 78691 174149 78716 174183
rect 78649 174141 78716 174149
rect 101149 174183 101199 174191
rect 101149 174149 101157 174183
rect 101191 174149 101199 174183
rect 101149 174141 101199 174149
rect 123649 174183 123866 174191
rect 123649 174149 123657 174183
rect 123860 174149 123866 174183
rect 123649 174141 123866 174149
rect 146149 174183 146566 174191
rect 146149 174149 146157 174183
rect 146149 174148 146178 174149
rect 146552 174148 146566 174183
rect 146149 174141 146566 174148
rect 56156 174116 56191 174141
rect 78666 174116 78716 174141
rect 101166 174116 101266 174141
rect 123666 174116 123866 174141
rect 146166 174116 146566 174141
rect 56156 174034 56191 174052
rect 78666 174032 78716 174052
rect 101166 174035 101266 174052
rect 123666 174036 123866 174052
rect 146166 174033 146566 174052
rect 56139 151183 56199 151191
rect 56139 151149 56147 151183
rect 56191 151149 56199 151183
rect 56139 151141 56199 151149
rect 78649 151183 78716 151191
rect 78649 151149 78657 151183
rect 78691 151149 78716 151183
rect 78649 151141 78716 151149
rect 101149 151183 101199 151191
rect 101149 151149 101157 151183
rect 101191 151149 101199 151183
rect 101149 151141 101199 151149
rect 123649 151183 123866 151191
rect 123649 151149 123657 151183
rect 123860 151149 123866 151183
rect 123649 151141 123866 151149
rect 146149 151183 146566 151191
rect 146149 151149 146157 151183
rect 146149 151148 146178 151149
rect 146552 151148 146566 151183
rect 146149 151141 146566 151148
rect 56156 151116 56191 151141
rect 78666 151116 78716 151141
rect 101166 151116 101266 151141
rect 123666 151116 123866 151141
rect 146166 151116 146566 151141
rect 56156 151018 56191 151032
rect 78666 151015 78716 151032
rect 101166 151018 101266 151032
rect 123666 151006 123866 151032
rect 146166 151002 146566 151032
rect 56139 128183 56199 128191
rect 56139 128149 56147 128183
rect 56191 128149 56199 128183
rect 56139 128141 56199 128149
rect 78649 128183 78716 128191
rect 78649 128149 78657 128183
rect 78691 128149 78716 128183
rect 78649 128141 78716 128149
rect 101149 128183 101199 128191
rect 101149 128149 101157 128183
rect 101191 128149 101199 128183
rect 101149 128141 101199 128149
rect 123649 128183 123866 128191
rect 123649 128149 123657 128183
rect 123860 128149 123866 128183
rect 123649 128141 123866 128149
rect 146149 128183 146566 128191
rect 146149 128149 146157 128183
rect 146149 128148 146178 128149
rect 146552 128148 146566 128183
rect 146149 128141 146566 128148
rect 56156 128116 56191 128141
rect 78666 128116 78716 128141
rect 101166 128116 101266 128141
rect 123666 128116 123866 128141
rect 146166 128116 146566 128141
rect 56156 128000 56191 128016
rect 78666 127991 78716 128016
rect 101166 127995 101266 128016
rect 123666 127995 123866 128016
rect 146166 127984 146566 128016
rect 56139 105183 56199 105191
rect 56139 105149 56147 105183
rect 56191 105149 56199 105183
rect 56139 105141 56199 105149
rect 78649 105183 78716 105191
rect 78649 105149 78657 105183
rect 78691 105149 78716 105183
rect 78649 105141 78716 105149
rect 101149 105183 101199 105191
rect 101149 105149 101157 105183
rect 101191 105149 101199 105183
rect 101149 105141 101199 105149
rect 123649 105183 123866 105191
rect 123649 105149 123657 105183
rect 123860 105149 123866 105183
rect 123649 105141 123866 105149
rect 146149 105183 146566 105191
rect 146149 105149 146157 105183
rect 146149 105148 146178 105149
rect 146552 105148 146566 105183
rect 146149 105141 146566 105148
rect 56156 105116 56191 105141
rect 78666 105116 78716 105141
rect 101166 105116 101266 105141
rect 123666 105116 123866 105141
rect 146166 105116 146566 105141
rect 56156 104932 56191 104951
rect 78666 104931 78716 104951
rect 101166 104922 101266 104951
rect 123666 104917 123866 104951
rect 146166 104930 146566 104951
rect 56139 82183 56199 82191
rect 56139 82149 56147 82183
rect 56191 82149 56199 82183
rect 56139 82141 56199 82149
rect 78649 82183 78716 82191
rect 78649 82149 78657 82183
rect 78691 82149 78716 82183
rect 78649 82141 78716 82149
rect 101149 82183 101199 82191
rect 101149 82149 101157 82183
rect 101191 82149 101199 82183
rect 101149 82141 101199 82149
rect 123649 82183 123866 82191
rect 123649 82149 123657 82183
rect 123860 82149 123866 82183
rect 123649 82141 123866 82149
rect 146149 82183 146566 82191
rect 146149 82149 146157 82183
rect 146149 82148 146178 82149
rect 146552 82148 146566 82183
rect 146149 82141 146566 82148
rect 56156 82116 56191 82141
rect 78666 82116 78716 82141
rect 101166 82116 101266 82141
rect 123666 82116 123866 82141
rect 146166 82116 146566 82141
rect 56156 81801 56191 81816
rect 78666 81798 78716 81816
rect 101166 81789 101266 81816
rect 123666 81798 123866 81816
rect 146166 81794 146566 81816
rect 56139 59183 56199 59191
rect 56139 59149 56147 59183
rect 56191 59149 56199 59183
rect 56139 59141 56199 59149
rect 78649 59183 78716 59191
rect 78649 59149 78657 59183
rect 78691 59149 78716 59183
rect 78649 59141 78716 59149
rect 101149 59183 101199 59191
rect 101149 59149 101157 59183
rect 101191 59149 101199 59183
rect 101149 59141 101199 59149
rect 123649 59183 123866 59191
rect 123649 59149 123657 59183
rect 123860 59149 123866 59183
rect 123649 59141 123866 59149
rect 146149 59183 146566 59191
rect 146149 59149 146157 59183
rect 146149 59148 146178 59149
rect 146552 59148 146566 59183
rect 146149 59141 146566 59148
rect 56156 59116 56191 59141
rect 78666 59116 78716 59141
rect 101166 59116 101266 59141
rect 123666 59116 123866 59141
rect 146166 59116 146566 59141
rect 56156 58598 56191 58616
rect 78666 58594 78716 58616
rect 101166 58578 101266 58616
rect 123666 58578 123866 58616
rect 146166 58590 146566 58616
rect 56139 36183 56199 36191
rect 56139 36149 56147 36183
rect 56191 36149 56199 36183
rect 56139 36141 56199 36149
rect 78649 36183 78716 36191
rect 78649 36149 78657 36183
rect 78691 36149 78716 36183
rect 78649 36141 78716 36149
rect 101149 36183 101199 36191
rect 101149 36149 101157 36183
rect 101191 36149 101199 36183
rect 101149 36141 101199 36149
rect 123649 36183 123866 36191
rect 123649 36149 123657 36183
rect 123860 36149 123866 36183
rect 123649 36141 123866 36149
rect 146149 36183 146566 36191
rect 146149 36149 146157 36183
rect 146149 36148 146178 36149
rect 146552 36148 146566 36183
rect 146149 36141 146566 36148
rect 56156 36116 56191 36141
rect 78666 36116 78716 36141
rect 101166 36116 101266 36141
rect 123666 36116 123866 36141
rect 146166 36116 146566 36141
rect 56156 35388 56191 35416
rect 78666 35386 78716 35416
rect 101166 35393 101266 35416
rect 123666 35391 123866 35416
rect 146166 35395 146566 35416
rect 56139 13183 56199 13191
rect 56139 13149 56147 13183
rect 56191 13149 56199 13183
rect 56139 13141 56199 13149
rect 78649 13183 78716 13191
rect 78649 13149 78657 13183
rect 78691 13149 78716 13183
rect 78649 13141 78716 13149
rect 101149 13183 101199 13191
rect 101149 13149 101157 13183
rect 101191 13149 101199 13183
rect 101149 13141 101199 13149
rect 123649 13183 123866 13191
rect 123649 13149 123657 13183
rect 123860 13149 123866 13183
rect 123649 13141 123866 13149
rect 146149 13183 146566 13191
rect 146149 13149 146157 13183
rect 146149 13148 146178 13149
rect 146552 13148 146566 13183
rect 146149 13141 146566 13148
rect 56156 13116 56191 13141
rect 78666 13116 78716 13141
rect 101166 13116 101266 13141
rect 123666 13116 123866 13141
rect 146166 13116 146566 13141
rect 56156 3097 56191 3116
rect 78666 3084 78716 3116
rect 101166 3050 101266 3116
rect 123666 3058 123866 3116
rect 146166 3076 146566 3116
<< polycont >>
rect 56147 220149 56191 220183
rect 78657 220149 78691 220183
rect 101157 220149 101191 220183
rect 123657 220149 123860 220183
rect 146157 220149 146552 220183
rect 146178 220148 146552 220149
rect 56147 197149 56191 197183
rect 78657 197149 78691 197183
rect 101157 197149 101191 197183
rect 123657 197149 123860 197183
rect 146157 197149 146552 197183
rect 146178 197148 146552 197149
rect 56147 174149 56191 174183
rect 78657 174149 78691 174183
rect 101157 174149 101191 174183
rect 123657 174149 123860 174183
rect 146157 174149 146552 174183
rect 146178 174148 146552 174149
rect 56147 151149 56191 151183
rect 78657 151149 78691 151183
rect 101157 151149 101191 151183
rect 123657 151149 123860 151183
rect 146157 151149 146552 151183
rect 146178 151148 146552 151149
rect 56147 128149 56191 128183
rect 78657 128149 78691 128183
rect 101157 128149 101191 128183
rect 123657 128149 123860 128183
rect 146157 128149 146552 128183
rect 146178 128148 146552 128149
rect 56147 105149 56191 105183
rect 78657 105149 78691 105183
rect 101157 105149 101191 105183
rect 123657 105149 123860 105183
rect 146157 105149 146552 105183
rect 146178 105148 146552 105149
rect 56147 82149 56191 82183
rect 78657 82149 78691 82183
rect 101157 82149 101191 82183
rect 123657 82149 123860 82183
rect 146157 82149 146552 82183
rect 146178 82148 146552 82149
rect 56147 59149 56191 59183
rect 78657 59149 78691 59183
rect 101157 59149 101191 59183
rect 123657 59149 123860 59183
rect 146157 59149 146552 59183
rect 146178 59148 146552 59149
rect 56147 36149 56191 36183
rect 78657 36149 78691 36183
rect 101157 36149 101191 36183
rect 123657 36149 123860 36183
rect 146157 36149 146552 36183
rect 146178 36148 146552 36149
rect 56147 13149 56191 13183
rect 78657 13149 78691 13183
rect 101157 13149 101191 13183
rect 123657 13149 123860 13183
rect 146157 13149 146552 13183
rect 146178 13148 146552 13149
<< locali >>
rect 56139 220183 56199 220191
rect 56139 220149 56147 220183
rect 56191 220149 56199 220183
rect 56139 220141 56199 220149
rect 78649 220183 78716 220191
rect 78649 220149 78657 220183
rect 78691 220149 78716 220183
rect 78649 220141 78716 220149
rect 101149 220183 101199 220191
rect 101149 220149 101157 220183
rect 101191 220149 101199 220183
rect 101149 220141 101199 220149
rect 123649 220183 123866 220191
rect 123649 220149 123657 220183
rect 123860 220149 123866 220183
rect 123649 220141 123866 220149
rect 146149 220183 146566 220191
rect 146149 220149 146157 220183
rect 146149 220148 146178 220149
rect 146552 220148 146566 220183
rect 146149 220141 146566 220148
rect 55958 220103 56046 220114
rect 55958 220086 55964 220103
rect 56045 220086 56046 220103
rect 55958 220076 56046 220086
rect 56066 220103 56154 220114
rect 56066 220086 56068 220103
rect 56144 220086 56154 220103
rect 56066 220076 56154 220086
rect 56193 220103 56289 220114
rect 56193 220086 56203 220103
rect 56284 220086 56289 220103
rect 56193 220076 56289 220086
rect 78468 220103 78556 220114
rect 78468 220086 78474 220103
rect 78555 220086 78556 220103
rect 78468 220076 78556 220086
rect 78576 220103 78664 220114
rect 78576 220086 78578 220103
rect 78654 220086 78664 220103
rect 78576 220076 78664 220086
rect 78718 220103 78814 220114
rect 78718 220086 78728 220103
rect 78809 220086 78814 220103
rect 78718 220076 78814 220086
rect 100968 220103 101056 220114
rect 100968 220086 100974 220103
rect 101055 220086 101056 220103
rect 100968 220076 101056 220086
rect 101076 220103 101164 220114
rect 101076 220086 101078 220103
rect 101154 220086 101164 220103
rect 101076 220076 101164 220086
rect 101268 220103 101364 220114
rect 101268 220086 101278 220103
rect 101359 220086 101364 220103
rect 101268 220076 101364 220086
rect 123468 220103 123556 220114
rect 123468 220086 123474 220103
rect 123555 220086 123556 220103
rect 123468 220076 123556 220086
rect 123576 220103 123664 220114
rect 123576 220086 123578 220103
rect 123654 220086 123664 220103
rect 123576 220076 123664 220086
rect 123868 220103 123964 220114
rect 123868 220086 123878 220103
rect 123959 220086 123964 220103
rect 123868 220076 123964 220086
rect 145968 220103 146056 220114
rect 145968 220086 145974 220103
rect 146055 220086 146056 220103
rect 145968 220076 146056 220086
rect 146076 220103 146164 220114
rect 146076 220086 146078 220103
rect 146154 220086 146164 220103
rect 146076 220076 146164 220086
rect 146568 220103 146664 220114
rect 146568 220086 146578 220103
rect 146659 220086 146664 220103
rect 146568 220076 146664 220086
rect 56139 197183 56199 197191
rect 56139 197149 56147 197183
rect 56191 197149 56199 197183
rect 56139 197141 56199 197149
rect 78649 197183 78716 197191
rect 78649 197149 78657 197183
rect 78691 197149 78716 197183
rect 78649 197141 78716 197149
rect 101149 197183 101199 197191
rect 101149 197149 101157 197183
rect 101191 197149 101199 197183
rect 101149 197141 101199 197149
rect 123649 197183 123866 197191
rect 123649 197149 123657 197183
rect 123860 197149 123866 197183
rect 123649 197141 123866 197149
rect 146149 197183 146566 197191
rect 146149 197149 146157 197183
rect 146149 197148 146178 197149
rect 146552 197148 146566 197183
rect 146149 197141 146566 197148
rect 55958 197103 56046 197114
rect 55958 197073 55964 197103
rect 56045 197073 56046 197103
rect 55958 197063 56046 197073
rect 56066 197103 56154 197114
rect 56066 197073 56068 197103
rect 56144 197073 56154 197103
rect 56066 197063 56154 197073
rect 56193 197103 56289 197114
rect 56193 197073 56203 197103
rect 56284 197073 56289 197103
rect 56193 197063 56289 197073
rect 78468 197103 78556 197114
rect 78468 197073 78474 197103
rect 78555 197073 78556 197103
rect 78468 197063 78556 197073
rect 78576 197103 78664 197114
rect 78576 197073 78578 197103
rect 78654 197073 78664 197103
rect 78576 197063 78664 197073
rect 78718 197103 78814 197114
rect 78718 197073 78728 197103
rect 78809 197073 78814 197103
rect 78718 197063 78814 197073
rect 100968 197103 101056 197114
rect 100968 197073 100974 197103
rect 101055 197073 101056 197103
rect 100968 197063 101056 197073
rect 101076 197103 101164 197114
rect 101076 197073 101078 197103
rect 101154 197073 101164 197103
rect 101076 197063 101164 197073
rect 101268 197103 101364 197114
rect 101268 197073 101278 197103
rect 101359 197073 101364 197103
rect 101268 197063 101364 197073
rect 123468 197103 123556 197114
rect 123468 197073 123474 197103
rect 123555 197073 123556 197103
rect 123468 197063 123556 197073
rect 123576 197103 123664 197114
rect 123576 197073 123578 197103
rect 123654 197073 123664 197103
rect 123576 197063 123664 197073
rect 123868 197103 123964 197114
rect 123868 197073 123878 197103
rect 123959 197073 123964 197103
rect 123868 197063 123964 197073
rect 145968 197103 146056 197114
rect 145968 197073 145974 197103
rect 146055 197073 146056 197103
rect 145968 197063 146056 197073
rect 146076 197103 146164 197114
rect 146076 197073 146078 197103
rect 146154 197073 146164 197103
rect 146076 197063 146164 197073
rect 146568 197103 146664 197114
rect 146568 197073 146578 197103
rect 146659 197073 146664 197103
rect 146568 197063 146664 197073
rect 56139 174183 56199 174191
rect 56139 174149 56147 174183
rect 56191 174149 56199 174183
rect 56139 174141 56199 174149
rect 78649 174183 78716 174191
rect 78649 174149 78657 174183
rect 78691 174149 78716 174183
rect 78649 174141 78716 174149
rect 101149 174183 101199 174191
rect 101149 174149 101157 174183
rect 101191 174149 101199 174183
rect 101149 174141 101199 174149
rect 123649 174183 123866 174191
rect 123649 174149 123657 174183
rect 123860 174149 123866 174183
rect 123649 174141 123866 174149
rect 146149 174183 146566 174191
rect 146149 174149 146157 174183
rect 146149 174148 146178 174149
rect 146552 174148 146566 174183
rect 146149 174141 146566 174148
rect 55958 174103 56046 174114
rect 55958 174064 55964 174103
rect 56045 174064 56046 174103
rect 55958 174054 56046 174064
rect 56066 174103 56154 174114
rect 56066 174064 56068 174103
rect 56144 174064 56154 174103
rect 56066 174054 56154 174064
rect 56193 174103 56289 174114
rect 56193 174064 56203 174103
rect 56284 174064 56289 174103
rect 56193 174054 56289 174064
rect 78468 174103 78556 174114
rect 78468 174064 78474 174103
rect 78555 174064 78556 174103
rect 78468 174054 78556 174064
rect 78576 174103 78664 174114
rect 78576 174064 78578 174103
rect 78654 174064 78664 174103
rect 78576 174054 78664 174064
rect 78718 174103 78814 174114
rect 78718 174064 78728 174103
rect 78809 174064 78814 174103
rect 78718 174054 78814 174064
rect 100968 174103 101056 174114
rect 100968 174064 100974 174103
rect 101055 174064 101056 174103
rect 100968 174054 101056 174064
rect 101076 174103 101164 174114
rect 101076 174064 101078 174103
rect 101154 174064 101164 174103
rect 101076 174054 101164 174064
rect 101268 174103 101364 174114
rect 101268 174064 101278 174103
rect 101359 174064 101364 174103
rect 101268 174054 101364 174064
rect 123468 174103 123556 174114
rect 123468 174064 123474 174103
rect 123555 174064 123556 174103
rect 123468 174054 123556 174064
rect 123576 174103 123664 174114
rect 123576 174064 123578 174103
rect 123654 174064 123664 174103
rect 123576 174054 123664 174064
rect 123868 174103 123964 174114
rect 123868 174064 123878 174103
rect 123959 174064 123964 174103
rect 123868 174054 123964 174064
rect 145968 174103 146056 174114
rect 145968 174064 145974 174103
rect 146055 174064 146056 174103
rect 145968 174054 146056 174064
rect 146076 174103 146164 174114
rect 146076 174064 146078 174103
rect 146154 174064 146164 174103
rect 146076 174054 146164 174064
rect 146568 174103 146664 174114
rect 146568 174064 146578 174103
rect 146659 174064 146664 174103
rect 146568 174054 146664 174064
rect 56139 151183 56199 151191
rect 56139 151149 56147 151183
rect 56191 151149 56199 151183
rect 56139 151141 56199 151149
rect 78649 151183 78716 151191
rect 78649 151149 78657 151183
rect 78691 151149 78716 151183
rect 78649 151141 78716 151149
rect 101149 151183 101199 151191
rect 101149 151149 101157 151183
rect 101191 151149 101199 151183
rect 101149 151141 101199 151149
rect 123649 151183 123866 151191
rect 123649 151149 123657 151183
rect 123860 151149 123866 151183
rect 123649 151141 123866 151149
rect 146149 151183 146566 151191
rect 146149 151149 146157 151183
rect 146149 151148 146178 151149
rect 146552 151148 146566 151183
rect 146149 151141 146566 151148
rect 55958 151103 56046 151114
rect 55958 151044 55964 151103
rect 56045 151044 56046 151103
rect 55958 151034 56046 151044
rect 56066 151103 56154 151114
rect 56066 151044 56068 151103
rect 56144 151044 56154 151103
rect 56066 151034 56154 151044
rect 56193 151103 56289 151114
rect 56193 151044 56203 151103
rect 56284 151044 56289 151103
rect 56193 151034 56289 151044
rect 78468 151103 78556 151114
rect 78468 151044 78474 151103
rect 78555 151044 78556 151103
rect 78468 151034 78556 151044
rect 78576 151103 78664 151114
rect 78576 151044 78578 151103
rect 78654 151044 78664 151103
rect 78576 151034 78664 151044
rect 78718 151103 78814 151114
rect 78718 151044 78728 151103
rect 78809 151044 78814 151103
rect 78718 151034 78814 151044
rect 100968 151103 101056 151114
rect 100968 151044 100974 151103
rect 101055 151044 101056 151103
rect 100968 151034 101056 151044
rect 101076 151103 101164 151114
rect 101076 151044 101078 151103
rect 101154 151044 101164 151103
rect 101076 151034 101164 151044
rect 101268 151103 101364 151114
rect 101268 151044 101278 151103
rect 101359 151044 101364 151103
rect 101268 151034 101364 151044
rect 123468 151103 123556 151114
rect 123468 151044 123474 151103
rect 123555 151044 123556 151103
rect 123468 151034 123556 151044
rect 123576 151103 123664 151114
rect 123576 151044 123578 151103
rect 123654 151044 123664 151103
rect 123576 151034 123664 151044
rect 123868 151103 123964 151114
rect 123868 151044 123878 151103
rect 123959 151044 123964 151103
rect 123868 151034 123964 151044
rect 145968 151103 146056 151114
rect 145968 151044 145974 151103
rect 146055 151044 146056 151103
rect 145968 151034 146056 151044
rect 146076 151103 146164 151114
rect 146076 151044 146078 151103
rect 146154 151044 146164 151103
rect 146076 151034 146164 151044
rect 146568 151103 146664 151114
rect 146568 151044 146578 151103
rect 146659 151044 146664 151103
rect 146568 151034 146664 151044
rect 56139 128183 56199 128191
rect 56139 128149 56147 128183
rect 56191 128149 56199 128183
rect 56139 128141 56199 128149
rect 78649 128183 78716 128191
rect 78649 128149 78657 128183
rect 78691 128149 78716 128183
rect 78649 128141 78716 128149
rect 101149 128183 101199 128191
rect 101149 128149 101157 128183
rect 101191 128149 101199 128183
rect 101149 128141 101199 128149
rect 123649 128183 123866 128191
rect 123649 128149 123657 128183
rect 123860 128149 123866 128183
rect 123649 128141 123866 128149
rect 146149 128183 146566 128191
rect 146149 128149 146157 128183
rect 146149 128148 146178 128149
rect 146552 128148 146566 128183
rect 146149 128141 146566 128148
rect 55958 128103 56046 128114
rect 55958 128028 55964 128103
rect 56045 128028 56046 128103
rect 55958 128018 56046 128028
rect 56066 128103 56154 128114
rect 56066 128028 56068 128103
rect 56144 128028 56154 128103
rect 56066 128018 56154 128028
rect 56193 128103 56289 128114
rect 56193 128028 56203 128103
rect 56284 128028 56289 128103
rect 56193 128018 56289 128028
rect 78468 128103 78556 128114
rect 78468 128028 78474 128103
rect 78555 128028 78556 128103
rect 78468 128018 78556 128028
rect 78576 128103 78664 128114
rect 78576 128028 78578 128103
rect 78654 128028 78664 128103
rect 78576 128018 78664 128028
rect 78718 128103 78814 128114
rect 78718 128028 78728 128103
rect 78809 128028 78814 128103
rect 78718 128018 78814 128028
rect 100968 128103 101056 128114
rect 100968 128028 100974 128103
rect 101055 128028 101056 128103
rect 100968 128018 101056 128028
rect 101076 128103 101164 128114
rect 101076 128028 101078 128103
rect 101154 128028 101164 128103
rect 101076 128018 101164 128028
rect 101268 128103 101364 128114
rect 101268 128028 101278 128103
rect 101359 128028 101364 128103
rect 101268 128018 101364 128028
rect 123468 128103 123556 128114
rect 123468 128028 123474 128103
rect 123555 128028 123556 128103
rect 123468 128018 123556 128028
rect 123576 128103 123664 128114
rect 123576 128028 123578 128103
rect 123654 128028 123664 128103
rect 123576 128018 123664 128028
rect 123868 128103 123964 128114
rect 123868 128028 123878 128103
rect 123959 128028 123964 128103
rect 123868 128018 123964 128028
rect 145968 128103 146056 128114
rect 145968 128028 145974 128103
rect 146055 128028 146056 128103
rect 145968 128018 146056 128028
rect 146076 128103 146164 128114
rect 146076 128028 146078 128103
rect 146154 128028 146164 128103
rect 146076 128018 146164 128028
rect 146568 128103 146664 128114
rect 146568 128028 146578 128103
rect 146659 128028 146664 128103
rect 146568 128018 146664 128028
rect 56139 105183 56199 105191
rect 56139 105149 56147 105183
rect 56191 105149 56199 105183
rect 56139 105141 56199 105149
rect 78649 105183 78716 105191
rect 78649 105149 78657 105183
rect 78691 105149 78716 105183
rect 78649 105141 78716 105149
rect 101149 105183 101199 105191
rect 101149 105149 101157 105183
rect 101191 105149 101199 105183
rect 101149 105141 101199 105149
rect 123649 105183 123866 105191
rect 123649 105149 123657 105183
rect 123860 105149 123866 105183
rect 123649 105141 123866 105149
rect 146149 105183 146566 105191
rect 146149 105149 146157 105183
rect 146149 105148 146178 105149
rect 146552 105148 146566 105183
rect 146149 105141 146566 105148
rect 55958 105103 56046 105114
rect 55958 104963 55964 105103
rect 56045 104963 56046 105103
rect 55958 104953 56046 104963
rect 56066 105103 56154 105114
rect 56066 104963 56068 105103
rect 56144 104963 56154 105103
rect 56066 104953 56154 104963
rect 56193 105103 56289 105114
rect 56193 104963 56203 105103
rect 56284 104963 56289 105103
rect 56193 104953 56289 104963
rect 78468 105103 78556 105114
rect 78468 104963 78474 105103
rect 78555 104963 78556 105103
rect 78468 104953 78556 104963
rect 78576 105103 78664 105114
rect 78576 104963 78578 105103
rect 78654 104963 78664 105103
rect 78576 104953 78664 104963
rect 78718 105103 78814 105114
rect 78718 104963 78728 105103
rect 78809 104963 78814 105103
rect 78718 104953 78814 104963
rect 100968 105103 101056 105114
rect 100968 104963 100974 105103
rect 101055 104963 101056 105103
rect 100968 104953 101056 104963
rect 101076 105103 101164 105114
rect 101076 104963 101078 105103
rect 101154 104963 101164 105103
rect 101076 104953 101164 104963
rect 101268 105103 101364 105114
rect 101268 104963 101278 105103
rect 101359 104963 101364 105103
rect 101268 104953 101364 104963
rect 123468 105103 123556 105114
rect 123468 104963 123474 105103
rect 123555 104963 123556 105103
rect 123468 104953 123556 104963
rect 123576 105103 123664 105114
rect 123576 104963 123578 105103
rect 123654 104963 123664 105103
rect 123576 104953 123664 104963
rect 123868 105103 123964 105114
rect 123868 104963 123878 105103
rect 123959 104963 123964 105103
rect 123868 104953 123964 104963
rect 145968 105103 146056 105114
rect 145968 104963 145974 105103
rect 146055 104963 146056 105103
rect 145968 104953 146056 104963
rect 146076 105103 146164 105114
rect 146076 104963 146078 105103
rect 146154 104963 146164 105103
rect 146076 104953 146164 104963
rect 146568 105103 146664 105114
rect 146568 104963 146578 105103
rect 146659 104963 146664 105103
rect 146568 104953 146664 104963
rect 56139 82183 56199 82191
rect 56139 82149 56147 82183
rect 56191 82149 56199 82183
rect 56139 82141 56199 82149
rect 78649 82183 78716 82191
rect 78649 82149 78657 82183
rect 78691 82149 78716 82183
rect 78649 82141 78716 82149
rect 101149 82183 101199 82191
rect 101149 82149 101157 82183
rect 101191 82149 101199 82183
rect 101149 82141 101199 82149
rect 123649 82183 123866 82191
rect 123649 82149 123657 82183
rect 123860 82149 123866 82183
rect 123649 82141 123866 82149
rect 146149 82183 146566 82191
rect 146149 82149 146157 82183
rect 146149 82148 146178 82149
rect 146552 82148 146566 82183
rect 146149 82141 146566 82148
rect 55958 82103 56046 82114
rect 55958 81828 55964 82103
rect 56045 81828 56046 82103
rect 55958 81818 56046 81828
rect 56066 82103 56154 82114
rect 56066 81828 56068 82103
rect 56144 81828 56154 82103
rect 56066 81818 56154 81828
rect 56193 82103 56289 82114
rect 56193 81828 56203 82103
rect 56284 81828 56289 82103
rect 56193 81818 56289 81828
rect 78468 82103 78556 82114
rect 78468 81828 78474 82103
rect 78555 81828 78556 82103
rect 78468 81818 78556 81828
rect 78576 82103 78664 82114
rect 78576 81828 78578 82103
rect 78654 81828 78664 82103
rect 78576 81818 78664 81828
rect 78718 82103 78814 82114
rect 78718 81828 78728 82103
rect 78809 81828 78814 82103
rect 78718 81818 78814 81828
rect 100968 82103 101056 82114
rect 100968 81828 100974 82103
rect 101055 81828 101056 82103
rect 100968 81818 101056 81828
rect 101076 82103 101164 82114
rect 101076 81828 101078 82103
rect 101154 81828 101164 82103
rect 101076 81818 101164 81828
rect 101268 82103 101364 82114
rect 101268 81828 101278 82103
rect 101359 81828 101364 82103
rect 101268 81818 101364 81828
rect 123468 82103 123556 82114
rect 123468 81828 123474 82103
rect 123555 81828 123556 82103
rect 123468 81818 123556 81828
rect 123576 82103 123664 82114
rect 123576 81828 123578 82103
rect 123654 81828 123664 82103
rect 123576 81818 123664 81828
rect 123868 82103 123964 82114
rect 123868 81828 123878 82103
rect 123959 81828 123964 82103
rect 123868 81818 123964 81828
rect 145968 82103 146056 82114
rect 145968 81828 145974 82103
rect 146055 81828 146056 82103
rect 145968 81818 146056 81828
rect 146076 82103 146164 82114
rect 146076 81828 146078 82103
rect 146154 81828 146164 82103
rect 146076 81818 146164 81828
rect 146568 82103 146664 82114
rect 146568 81828 146578 82103
rect 146659 81828 146664 82103
rect 146568 81818 146664 81828
rect 56139 59183 56199 59191
rect 56139 59149 56147 59183
rect 56191 59149 56199 59183
rect 56139 59141 56199 59149
rect 78649 59183 78716 59191
rect 78649 59149 78657 59183
rect 78691 59149 78716 59183
rect 78649 59141 78716 59149
rect 101149 59183 101199 59191
rect 101149 59149 101157 59183
rect 101191 59149 101199 59183
rect 101149 59141 101199 59149
rect 123649 59183 123866 59191
rect 123649 59149 123657 59183
rect 123860 59149 123866 59183
rect 123649 59141 123866 59149
rect 146149 59183 146566 59191
rect 146149 59149 146157 59183
rect 146149 59148 146178 59149
rect 146552 59148 146566 59183
rect 146149 59141 146566 59148
rect 55958 59103 56046 59114
rect 55958 58628 55964 59103
rect 56045 58628 56046 59103
rect 55958 58618 56046 58628
rect 56066 59103 56154 59114
rect 56066 58628 56068 59103
rect 56144 58628 56154 59103
rect 56066 58618 56154 58628
rect 56193 59103 56289 59114
rect 56193 58628 56203 59103
rect 56284 58628 56289 59103
rect 56193 58618 56289 58628
rect 78468 59103 78556 59114
rect 78468 58628 78474 59103
rect 78555 58628 78556 59103
rect 78468 58618 78556 58628
rect 78576 59103 78664 59114
rect 78576 58628 78578 59103
rect 78654 58628 78664 59103
rect 78576 58618 78664 58628
rect 78718 59103 78814 59114
rect 78718 58628 78728 59103
rect 78809 58628 78814 59103
rect 78718 58618 78814 58628
rect 100968 59103 101056 59114
rect 100968 58628 100974 59103
rect 101055 58628 101056 59103
rect 100968 58618 101056 58628
rect 101076 59103 101164 59114
rect 101076 58628 101078 59103
rect 101154 58628 101164 59103
rect 101076 58618 101164 58628
rect 101268 59103 101364 59114
rect 101268 58628 101278 59103
rect 101359 58628 101364 59103
rect 101268 58618 101364 58628
rect 123468 59103 123556 59114
rect 123468 58628 123474 59103
rect 123555 58628 123556 59103
rect 123468 58618 123556 58628
rect 123576 59103 123664 59114
rect 123576 58628 123578 59103
rect 123654 58628 123664 59103
rect 123576 58618 123664 58628
rect 123868 59103 123964 59114
rect 123868 58628 123878 59103
rect 123959 58628 123964 59103
rect 123868 58618 123964 58628
rect 145968 59103 146056 59114
rect 145968 58628 145974 59103
rect 146055 58628 146056 59103
rect 145968 58618 146056 58628
rect 146076 59103 146164 59114
rect 146076 58628 146078 59103
rect 146154 58628 146164 59103
rect 146076 58618 146164 58628
rect 146568 59103 146664 59114
rect 146568 58628 146578 59103
rect 146659 58628 146664 59103
rect 146568 58618 146664 58628
rect 56139 36183 56199 36191
rect 56139 36149 56147 36183
rect 56191 36149 56199 36183
rect 56139 36141 56199 36149
rect 78649 36183 78716 36191
rect 78649 36149 78657 36183
rect 78691 36149 78716 36183
rect 78649 36141 78716 36149
rect 101149 36183 101199 36191
rect 101149 36149 101157 36183
rect 101191 36149 101199 36183
rect 101149 36141 101199 36149
rect 123649 36183 123866 36191
rect 123649 36149 123657 36183
rect 123860 36149 123866 36183
rect 123649 36141 123866 36149
rect 146149 36183 146566 36191
rect 146149 36149 146157 36183
rect 146149 36148 146178 36149
rect 146552 36148 146566 36183
rect 146149 36141 146566 36148
rect 55958 36103 56046 36114
rect 55958 35428 55964 36103
rect 56045 35428 56046 36103
rect 55958 35418 56046 35428
rect 56066 36103 56154 36114
rect 56066 35428 56068 36103
rect 56144 35428 56154 36103
rect 56066 35418 56154 35428
rect 56193 36103 56289 36114
rect 56193 35428 56203 36103
rect 56284 35428 56289 36103
rect 56193 35418 56289 35428
rect 78468 36103 78556 36114
rect 78468 35428 78474 36103
rect 78555 35428 78556 36103
rect 78468 35418 78556 35428
rect 78576 36103 78664 36114
rect 78576 35428 78578 36103
rect 78654 35428 78664 36103
rect 78576 35418 78664 35428
rect 78718 36103 78814 36114
rect 78718 35428 78728 36103
rect 78809 35428 78814 36103
rect 78718 35418 78814 35428
rect 100968 36103 101056 36114
rect 100968 35428 100974 36103
rect 101055 35428 101056 36103
rect 100968 35418 101056 35428
rect 101076 36103 101164 36114
rect 101076 35428 101078 36103
rect 101154 35428 101164 36103
rect 101076 35418 101164 35428
rect 101268 36103 101364 36114
rect 101268 35428 101278 36103
rect 101359 35428 101364 36103
rect 101268 35418 101364 35428
rect 123468 36103 123556 36114
rect 123468 35428 123474 36103
rect 123555 35428 123556 36103
rect 123468 35418 123556 35428
rect 123576 36103 123664 36114
rect 123576 35428 123578 36103
rect 123654 35428 123664 36103
rect 123576 35418 123664 35428
rect 123868 36103 123964 36114
rect 123868 35428 123878 36103
rect 123959 35428 123964 36103
rect 123868 35418 123964 35428
rect 145968 36103 146056 36114
rect 145968 35428 145974 36103
rect 146055 35428 146056 36103
rect 145968 35418 146056 35428
rect 146076 36103 146164 36114
rect 146076 35428 146078 36103
rect 146154 35428 146164 36103
rect 146076 35418 146164 35428
rect 146568 36103 146664 36114
rect 146568 35428 146578 36103
rect 146659 35428 146664 36103
rect 146568 35418 146664 35428
rect 56139 13183 56199 13191
rect 56139 13149 56147 13183
rect 56191 13149 56199 13183
rect 56139 13141 56199 13149
rect 78649 13183 78716 13191
rect 78649 13149 78657 13183
rect 78691 13149 78716 13183
rect 78649 13141 78716 13149
rect 101149 13183 101199 13191
rect 101149 13149 101157 13183
rect 101191 13149 101199 13183
rect 101149 13141 101199 13149
rect 123649 13183 123866 13191
rect 123649 13149 123657 13183
rect 123860 13149 123866 13183
rect 123649 13141 123866 13149
rect 146149 13183 146566 13191
rect 146149 13149 146157 13183
rect 146149 13148 146178 13149
rect 146552 13148 146566 13183
rect 146149 13141 146566 13148
rect 55958 13103 56046 13114
rect 55958 3128 55964 13103
rect 56045 3128 56046 13103
rect 55958 3118 56046 3128
rect 56066 13103 56154 13114
rect 56066 3128 56068 13103
rect 56144 3128 56154 13103
rect 56066 3118 56154 3128
rect 56193 13103 56289 13114
rect 56193 3128 56203 13103
rect 56284 3128 56289 13103
rect 56193 3118 56289 3128
rect 78468 13103 78556 13114
rect 78468 3128 78474 13103
rect 78555 3128 78556 13103
rect 78468 3118 78556 3128
rect 78576 13103 78664 13114
rect 78576 3128 78578 13103
rect 78654 3128 78664 13103
rect 78576 3118 78664 3128
rect 78718 13103 78814 13114
rect 78718 3128 78728 13103
rect 78809 3128 78814 13103
rect 78718 3118 78814 3128
rect 100968 13103 101056 13114
rect 100968 3128 100974 13103
rect 101055 3128 101056 13103
rect 100968 3118 101056 3128
rect 101076 13103 101164 13114
rect 101076 3128 101078 13103
rect 101154 3128 101164 13103
rect 101076 3118 101164 3128
rect 101268 13103 101364 13114
rect 101268 3128 101278 13103
rect 101359 3128 101364 13103
rect 101268 3118 101364 3128
rect 123468 13103 123556 13114
rect 123468 3128 123474 13103
rect 123555 3128 123556 13103
rect 123468 3118 123556 3128
rect 123576 13103 123664 13114
rect 123576 3128 123578 13103
rect 123654 3128 123664 13103
rect 123576 3118 123664 3128
rect 123868 13103 123964 13114
rect 123868 3128 123878 13103
rect 123959 3128 123964 13103
rect 123868 3118 123964 3128
rect 145968 13103 146056 13114
rect 145968 3128 145974 13103
rect 146055 3128 146056 13103
rect 145968 3118 146056 3128
rect 146076 13103 146164 13114
rect 146076 3128 146078 13103
rect 146154 3128 146164 13103
rect 146076 3118 146164 3128
rect 146568 13103 146664 13114
rect 146568 3128 146578 13103
rect 146659 3128 146664 13103
rect 146568 3118 146664 3128
<< viali >>
rect 56147 220150 56191 220183
rect 78657 220150 78691 220183
rect 101157 220150 101191 220183
rect 123657 220150 123860 220183
rect 123691 220149 123860 220150
rect 146157 220150 146552 220183
rect 146178 220148 146552 220150
rect 55964 220086 55969 220103
rect 55969 220086 56028 220103
rect 56073 220086 56137 220103
rect 56209 220086 56279 220103
rect 56279 220086 56284 220103
rect 78474 220086 78479 220103
rect 78479 220086 78538 220103
rect 78583 220086 78647 220103
rect 78734 220086 78804 220103
rect 78804 220086 78809 220103
rect 100974 220086 100979 220103
rect 100979 220086 101038 220103
rect 101083 220086 101147 220103
rect 101284 220086 101354 220103
rect 101354 220086 101359 220103
rect 123474 220086 123479 220103
rect 123479 220086 123538 220103
rect 123583 220086 123647 220103
rect 123884 220086 123954 220103
rect 123954 220086 123959 220103
rect 145974 220086 145979 220103
rect 145979 220086 146038 220103
rect 146083 220086 146147 220103
rect 146584 220086 146654 220103
rect 146654 220086 146659 220103
rect 56147 197150 56191 197183
rect 78657 197150 78691 197183
rect 101157 197150 101191 197183
rect 123657 197150 123860 197183
rect 123691 197149 123860 197150
rect 146157 197150 146552 197183
rect 146178 197148 146552 197150
rect 55964 197073 55969 197103
rect 55969 197073 56028 197103
rect 56073 197073 56137 197103
rect 56209 197073 56279 197103
rect 56279 197073 56284 197103
rect 78474 197073 78479 197103
rect 78479 197073 78538 197103
rect 78583 197073 78647 197103
rect 78734 197073 78804 197103
rect 78804 197073 78809 197103
rect 100974 197073 100979 197103
rect 100979 197073 101038 197103
rect 101083 197073 101147 197103
rect 101284 197073 101354 197103
rect 101354 197073 101359 197103
rect 123474 197073 123479 197103
rect 123479 197073 123538 197103
rect 123583 197073 123647 197103
rect 123884 197073 123954 197103
rect 123954 197073 123959 197103
rect 145974 197073 145979 197103
rect 145979 197073 146038 197103
rect 146083 197073 146147 197103
rect 146584 197073 146654 197103
rect 146654 197073 146659 197103
rect 56147 174150 56191 174183
rect 78657 174150 78691 174183
rect 101157 174150 101191 174183
rect 123657 174150 123860 174183
rect 123691 174149 123860 174150
rect 146157 174150 146552 174183
rect 146178 174148 146552 174150
rect 55964 174064 55969 174103
rect 55969 174064 56028 174103
rect 56073 174064 56137 174103
rect 56209 174064 56279 174103
rect 56279 174064 56284 174103
rect 78474 174064 78479 174103
rect 78479 174064 78538 174103
rect 78583 174064 78647 174103
rect 78734 174064 78804 174103
rect 78804 174064 78809 174103
rect 100974 174064 100979 174103
rect 100979 174064 101038 174103
rect 101083 174064 101147 174103
rect 101284 174064 101354 174103
rect 101354 174064 101359 174103
rect 123474 174064 123479 174103
rect 123479 174064 123538 174103
rect 123583 174064 123647 174103
rect 123884 174064 123954 174103
rect 123954 174064 123959 174103
rect 145974 174064 145979 174103
rect 145979 174064 146038 174103
rect 146083 174064 146147 174103
rect 146584 174064 146654 174103
rect 146654 174064 146659 174103
rect 56147 151150 56191 151183
rect 78657 151150 78691 151183
rect 101157 151150 101191 151183
rect 123657 151150 123860 151183
rect 123691 151149 123860 151150
rect 146157 151150 146552 151183
rect 146178 151148 146552 151150
rect 55964 151044 55969 151103
rect 55969 151044 56028 151103
rect 56073 151044 56137 151103
rect 56209 151044 56279 151103
rect 56279 151044 56284 151103
rect 78474 151044 78479 151103
rect 78479 151044 78538 151103
rect 78583 151044 78647 151103
rect 78734 151044 78804 151103
rect 78804 151044 78809 151103
rect 100974 151044 100979 151103
rect 100979 151044 101038 151103
rect 101083 151044 101147 151103
rect 101284 151044 101354 151103
rect 101354 151044 101359 151103
rect 123474 151044 123479 151103
rect 123479 151044 123538 151103
rect 123583 151044 123647 151103
rect 123884 151044 123954 151103
rect 123954 151044 123959 151103
rect 145974 151044 145979 151103
rect 145979 151044 146038 151103
rect 146083 151044 146147 151103
rect 146584 151044 146654 151103
rect 146654 151044 146659 151103
rect 56147 128150 56191 128183
rect 78657 128150 78691 128183
rect 101157 128150 101191 128183
rect 123657 128150 123860 128183
rect 123691 128149 123860 128150
rect 146157 128150 146552 128183
rect 146178 128148 146552 128150
rect 55964 128028 55969 128103
rect 55969 128028 56028 128103
rect 56073 128028 56137 128103
rect 56209 128028 56279 128103
rect 56279 128028 56284 128103
rect 78474 128028 78479 128103
rect 78479 128028 78538 128103
rect 78583 128028 78647 128103
rect 78734 128028 78804 128103
rect 78804 128028 78809 128103
rect 100974 128028 100979 128103
rect 100979 128028 101038 128103
rect 101083 128028 101147 128103
rect 101284 128028 101354 128103
rect 101354 128028 101359 128103
rect 123474 128028 123479 128103
rect 123479 128028 123538 128103
rect 123583 128028 123647 128103
rect 123884 128028 123954 128103
rect 123954 128028 123959 128103
rect 145974 128028 145979 128103
rect 145979 128028 146038 128103
rect 146083 128028 146147 128103
rect 146584 128028 146654 128103
rect 146654 128028 146659 128103
rect 56147 105150 56191 105183
rect 78657 105150 78691 105183
rect 101157 105150 101191 105183
rect 123657 105150 123860 105183
rect 123691 105149 123860 105150
rect 146157 105150 146552 105183
rect 146178 105148 146552 105150
rect 55964 104963 55969 105103
rect 55969 104963 56028 105103
rect 56073 104963 56137 105103
rect 56209 104963 56279 105103
rect 56279 104963 56284 105103
rect 78474 104963 78479 105103
rect 78479 104963 78538 105103
rect 78583 104963 78647 105103
rect 78734 104963 78804 105103
rect 78804 104963 78809 105103
rect 100974 104963 100979 105103
rect 100979 104963 101038 105103
rect 101083 104963 101147 105103
rect 101284 104963 101354 105103
rect 101354 104963 101359 105103
rect 123474 104963 123479 105103
rect 123479 104963 123538 105103
rect 123583 104963 123647 105103
rect 123884 104963 123954 105103
rect 123954 104963 123959 105103
rect 145974 104963 145979 105103
rect 145979 104963 146038 105103
rect 146083 104963 146147 105103
rect 146584 104963 146654 105103
rect 146654 104963 146659 105103
rect 56147 82150 56191 82183
rect 78657 82150 78691 82183
rect 101157 82150 101191 82183
rect 123657 82150 123860 82183
rect 123691 82149 123860 82150
rect 146157 82150 146552 82183
rect 146178 82148 146552 82150
rect 55964 81828 55969 82103
rect 55969 81828 56028 82103
rect 56073 81828 56137 82103
rect 56209 81828 56279 82103
rect 56279 81828 56284 82103
rect 78474 81828 78479 82103
rect 78479 81828 78538 82103
rect 78583 81828 78647 82103
rect 78734 81828 78804 82103
rect 78804 81828 78809 82103
rect 100974 81828 100979 82103
rect 100979 81828 101038 82103
rect 101083 81828 101147 82103
rect 101284 81828 101354 82103
rect 101354 81828 101359 82103
rect 123474 81828 123479 82103
rect 123479 81828 123538 82103
rect 123583 81828 123647 82103
rect 123884 81828 123954 82103
rect 123954 81828 123959 82103
rect 145974 81828 145979 82103
rect 145979 81828 146038 82103
rect 146083 81828 146147 82103
rect 146584 81828 146654 82103
rect 146654 81828 146659 82103
rect 56147 59150 56191 59183
rect 78657 59150 78691 59183
rect 101157 59150 101191 59183
rect 123657 59150 123860 59183
rect 123691 59149 123860 59150
rect 146157 59150 146552 59183
rect 146178 59148 146552 59150
rect 55964 58628 55969 59103
rect 55969 58628 56028 59103
rect 56073 58628 56137 59103
rect 56209 58628 56279 59103
rect 56279 58628 56284 59103
rect 78474 58628 78479 59103
rect 78479 58628 78538 59103
rect 78583 58628 78647 59103
rect 78734 58628 78804 59103
rect 78804 58628 78809 59103
rect 100974 58628 100979 59103
rect 100979 58628 101038 59103
rect 101083 58628 101147 59103
rect 101284 58628 101354 59103
rect 101354 58628 101359 59103
rect 123474 58628 123479 59103
rect 123479 58628 123538 59103
rect 123583 58628 123647 59103
rect 123884 58628 123954 59103
rect 123954 58628 123959 59103
rect 145974 58628 145979 59103
rect 145979 58628 146038 59103
rect 146083 58628 146147 59103
rect 146584 58628 146654 59103
rect 146654 58628 146659 59103
rect 56147 36150 56191 36183
rect 78657 36150 78691 36183
rect 101157 36150 101191 36183
rect 123657 36150 123860 36183
rect 123691 36149 123860 36150
rect 146157 36150 146552 36183
rect 146178 36148 146552 36150
rect 55964 35428 55969 36103
rect 55969 35428 56028 36103
rect 56073 35428 56137 36103
rect 56209 35428 56279 36103
rect 56279 35428 56284 36103
rect 78474 35428 78479 36103
rect 78479 35428 78538 36103
rect 78583 35428 78647 36103
rect 78734 35428 78804 36103
rect 78804 35428 78809 36103
rect 100974 35428 100979 36103
rect 100979 35428 101038 36103
rect 101083 35428 101147 36103
rect 101284 35428 101354 36103
rect 101354 35428 101359 36103
rect 123474 35428 123479 36103
rect 123479 35428 123538 36103
rect 123583 35428 123647 36103
rect 123884 35428 123954 36103
rect 123954 35428 123959 36103
rect 145974 35428 145979 36103
rect 145979 35428 146038 36103
rect 146083 35428 146147 36103
rect 146584 35428 146654 36103
rect 146654 35428 146659 36103
rect 56147 13150 56191 13183
rect 78657 13150 78691 13183
rect 101157 13150 101191 13183
rect 123657 13150 123860 13183
rect 123691 13149 123860 13150
rect 146157 13150 146552 13183
rect 146178 13148 146552 13150
rect 55964 3128 55969 13103
rect 55969 3128 56028 13103
rect 56073 3128 56137 13103
rect 56209 3128 56279 13103
rect 56279 3128 56284 13103
rect 78474 3128 78479 13103
rect 78479 3128 78538 13103
rect 78583 3128 78647 13103
rect 78734 3128 78804 13103
rect 78804 3128 78809 13103
rect 100974 3128 100979 13103
rect 100979 3128 101038 13103
rect 101083 3128 101147 13103
rect 101284 3128 101354 13103
rect 101354 3128 101359 13103
rect 123474 3128 123479 13103
rect 123479 3128 123538 13103
rect 123583 3128 123647 13103
rect 123884 3128 123954 13103
rect 123954 3128 123959 13103
rect 145974 3128 145979 13103
rect 145979 3128 146038 13103
rect 146083 3128 146147 13103
rect 146584 3128 146654 13103
rect 146654 3128 146659 13103
<< metal1 >>
rect 54745 220515 56245 221020
rect 77245 220515 78745 221020
rect 99745 220515 101245 221020
rect 122245 220515 123745 221020
rect 144745 220515 146245 221020
rect 55958 220307 56035 220515
rect 78468 220307 78545 220515
rect 100968 220307 101045 220515
rect 123468 220307 123545 220515
rect 145968 220307 146045 220515
rect 55958 220103 56036 220307
rect 57750 220203 58024 220204
rect 56139 220183 58024 220203
rect 56139 220150 56147 220183
rect 56191 220150 58024 220183
rect 56139 220141 58024 220150
rect 55958 220086 55964 220103
rect 56028 220086 56036 220103
rect 55958 220077 56036 220086
rect 56066 220103 56144 220113
rect 56066 220086 56073 220103
rect 56137 220086 56144 220103
rect 56066 219916 56144 220086
rect 56065 219896 56144 219916
rect 56203 220103 56291 220114
rect 56203 220086 56209 220103
rect 56284 220086 56291 220103
rect 56203 220071 56291 220086
rect 78468 220103 78546 220307
rect 78649 220183 80532 220203
rect 78649 220150 78657 220183
rect 78691 220150 80532 220183
rect 78649 220141 80532 220150
rect 78468 220086 78474 220103
rect 78538 220086 78546 220103
rect 78468 220077 78546 220086
rect 78576 220103 78654 220113
rect 78576 220086 78583 220103
rect 78647 220086 78654 220103
rect 56065 219839 56143 219896
rect 55873 219771 56143 219839
rect 56203 219853 56281 220071
rect 78576 219916 78654 220086
rect 78575 219896 78654 219916
rect 78728 220103 78816 220114
rect 78728 220086 78734 220103
rect 78809 220086 78816 220103
rect 78728 220071 78816 220086
rect 100968 220103 101046 220307
rect 101149 220183 103018 220203
rect 101149 220150 101157 220183
rect 101191 220150 103018 220183
rect 101149 220141 103018 220150
rect 100968 220086 100974 220103
rect 101038 220086 101046 220103
rect 100968 220077 101046 220086
rect 101076 220103 101154 220113
rect 101076 220086 101083 220103
rect 101147 220086 101154 220103
rect 56203 219802 56691 219853
rect 78575 219839 78653 219896
rect 55873 219763 56142 219771
rect 55208 219762 56142 219763
rect 53983 219755 54481 219761
rect 54745 219755 56142 219762
rect 53983 219728 56142 219755
rect 56204 219733 56691 219802
rect 78373 219771 78653 219839
rect 78728 219853 78806 220071
rect 101076 219916 101154 220086
rect 101278 220103 101366 220114
rect 101278 220086 101284 220103
rect 101359 220086 101366 220103
rect 101278 220071 101366 220086
rect 123468 220103 123546 220307
rect 123649 220183 125532 220203
rect 123649 220150 123657 220183
rect 123649 220149 123691 220150
rect 123860 220149 125532 220183
rect 123649 220141 125532 220149
rect 125242 220140 125532 220141
rect 123468 220086 123474 220103
rect 123538 220086 123546 220103
rect 123468 220077 123546 220086
rect 123576 220103 123654 220113
rect 123576 220086 123583 220103
rect 123647 220086 123654 220103
rect 101278 220031 101356 220071
rect 101075 219896 101154 219916
rect 78728 219802 79191 219853
rect 101075 219839 101153 219896
rect 101277 219853 101357 220031
rect 123576 219916 123654 220086
rect 123575 219896 123654 219916
rect 123878 220103 123966 220114
rect 123878 220086 123884 220103
rect 123959 220098 123966 220103
rect 145968 220103 146046 220307
rect 146149 220183 148021 220203
rect 146149 220150 146157 220183
rect 146149 220148 146178 220150
rect 146552 220148 148021 220183
rect 146149 220141 148021 220148
rect 123959 220086 123971 220098
rect 53983 219327 55939 219728
rect 56064 219725 56142 219728
rect 56225 219626 56691 219733
rect 53983 218470 54481 219327
rect 54745 219321 55939 219327
rect 54745 219319 55224 219321
rect 53915 217940 54620 218470
rect 56256 216767 56691 219626
rect 76480 219761 76989 219764
rect 78373 219763 78652 219771
rect 77708 219762 78652 219763
rect 77245 219761 78652 219762
rect 76480 219728 78652 219761
rect 78729 219733 79191 219802
rect 100873 219771 101153 219839
rect 100873 219763 101152 219771
rect 100208 219762 101152 219763
rect 99745 219760 101152 219762
rect 99230 219750 101152 219760
rect 76480 219321 78449 219728
rect 78574 219725 78652 219728
rect 76480 219320 77724 219321
rect 76480 218560 76989 219320
rect 77245 219319 77724 219320
rect 76335 217850 77175 218560
rect 78756 216815 79191 219733
rect 98977 219728 101152 219750
rect 101273 219732 101691 219853
rect 123575 219839 123653 219896
rect 123878 219853 123971 220086
rect 145968 220086 145974 220103
rect 146038 220086 146046 220103
rect 145968 220077 146046 220086
rect 146076 220103 146154 220113
rect 146076 220086 146083 220103
rect 146147 220086 146154 220103
rect 146076 219916 146154 220086
rect 146578 220103 146666 220114
rect 146578 220086 146584 220103
rect 146659 220086 146666 220103
rect 146578 220081 146666 220086
rect 146075 219896 146154 219916
rect 123373 219771 123653 219839
rect 123373 219763 123652 219771
rect 122708 219762 123652 219763
rect 98977 219321 100949 219728
rect 101074 219725 101152 219728
rect 98977 218665 99481 219321
rect 99745 219319 100224 219321
rect 98865 217955 99705 218665
rect 101256 216843 101691 219732
rect 121480 219728 123652 219762
rect 121480 219321 123449 219728
rect 123574 219725 123652 219728
rect 121480 219320 122724 219321
rect 121480 218815 121960 219320
rect 122245 219319 122724 219320
rect 121400 217885 122000 218815
rect 123756 216846 124191 219853
rect 146075 219839 146153 219896
rect 146577 219853 146667 220081
rect 145873 219771 146153 219839
rect 145873 219763 146152 219771
rect 145208 219762 146152 219763
rect 143980 219728 146152 219762
rect 143980 219321 145949 219728
rect 146074 219725 146152 219728
rect 143980 219319 145224 219321
rect 143980 219318 144920 219319
rect 143980 218860 144484 219318
rect 143920 217930 144520 218860
rect 146256 216975 146691 219853
rect 56240 216330 56696 216767
rect 78744 216612 79191 216815
rect 78744 216452 79192 216612
rect 101246 216602 101691 216843
rect 78744 216374 79179 216452
rect 101246 216218 101690 216602
rect 123738 216293 124200 216846
rect 146150 216045 146750 216975
rect 55798 197325 56242 197641
rect 55958 197103 56036 197325
rect 58010 197204 58515 197368
rect 78407 197351 78609 197561
rect 57750 197203 58515 197204
rect 56139 197183 58515 197203
rect 56139 197150 56147 197183
rect 56191 197150 58515 197183
rect 56139 197141 58515 197150
rect 55958 197073 55964 197103
rect 56028 197073 56036 197103
rect 55958 197064 56036 197073
rect 56066 197103 56144 197113
rect 56066 197073 56073 197103
rect 56137 197073 56144 197103
rect 56066 196916 56144 197073
rect 56065 196896 56144 196916
rect 56203 197103 56291 197114
rect 56203 197073 56209 197103
rect 56284 197073 56291 197103
rect 56203 197061 56291 197073
rect 56065 196839 56143 196896
rect 55873 196771 56143 196839
rect 56203 196853 56281 197061
rect 56203 196802 56691 196853
rect 55873 196763 56142 196771
rect 55208 196762 56142 196763
rect 53983 196755 54481 196761
rect 54745 196755 56142 196762
rect 53983 196728 56142 196755
rect 56204 196733 56691 196802
rect 53983 196327 55939 196728
rect 56064 196725 56142 196728
rect 56225 196626 56691 196733
rect 53983 195250 54481 196327
rect 54745 196321 55939 196327
rect 54745 196319 55224 196321
rect 53980 193650 54485 195250
rect 56256 193985 56691 196626
rect 58010 195755 58515 197141
rect 78468 197307 78545 197351
rect 78468 197103 78546 197307
rect 80510 197203 81015 197368
rect 100788 197356 101240 197866
rect 78649 197183 81015 197203
rect 78649 197150 78657 197183
rect 78691 197150 81015 197183
rect 78649 197141 81015 197150
rect 78468 197073 78474 197103
rect 78538 197073 78546 197103
rect 78468 197064 78546 197073
rect 78576 197103 78654 197113
rect 78576 197073 78583 197103
rect 78647 197073 78654 197103
rect 78576 196916 78654 197073
rect 78575 196896 78654 196916
rect 78728 197103 78816 197114
rect 78728 197073 78734 197103
rect 78809 197073 78816 197103
rect 78728 197061 78816 197073
rect 78575 196839 78653 196896
rect 78373 196771 78653 196839
rect 78728 196853 78806 197061
rect 78728 196802 79191 196853
rect 76480 196761 76989 196764
rect 78373 196763 78652 196771
rect 77708 196762 78652 196763
rect 77245 196761 78652 196762
rect 76480 196728 78652 196761
rect 78729 196733 79191 196802
rect 76480 196321 78449 196728
rect 78574 196725 78652 196728
rect 76480 196320 77724 196321
rect 76480 195242 76989 196320
rect 77245 196319 77724 196320
rect 56200 192750 56970 193985
rect 76480 193650 76985 195242
rect 78756 193850 79191 196733
rect 80510 195755 81015 197141
rect 100968 197307 101045 197356
rect 100968 197103 101046 197307
rect 103010 197203 103515 197368
rect 123259 197361 123733 197793
rect 101149 197183 103515 197203
rect 101149 197150 101157 197183
rect 101191 197150 103515 197183
rect 101149 197141 103515 197150
rect 100968 197073 100974 197103
rect 101038 197073 101046 197103
rect 100968 197064 101046 197073
rect 101076 197103 101154 197113
rect 101076 197073 101083 197103
rect 101147 197073 101154 197103
rect 101076 196916 101154 197073
rect 101278 197103 101366 197114
rect 101278 197073 101284 197103
rect 101359 197073 101366 197103
rect 101278 197061 101366 197073
rect 101278 197031 101356 197061
rect 101075 196896 101154 196916
rect 101075 196839 101153 196896
rect 101277 196853 101357 197031
rect 100873 196771 101153 196839
rect 100873 196763 101152 196771
rect 100208 196762 101152 196763
rect 99745 196760 101152 196762
rect 99230 196750 101152 196760
rect 98977 196728 101152 196750
rect 101273 196732 101691 196853
rect 98977 196321 100949 196728
rect 101074 196725 101152 196728
rect 98977 195250 99481 196321
rect 99745 196319 100224 196321
rect 98977 195223 99485 195250
rect 78495 192615 79265 193850
rect 98980 193650 99485 195223
rect 101256 193843 101691 196732
rect 103010 195755 103515 197141
rect 123468 197307 123545 197361
rect 123468 197103 123546 197307
rect 125510 197203 126015 197368
rect 145793 197353 146245 197801
rect 123649 197183 126015 197203
rect 123649 197150 123657 197183
rect 123649 197149 123691 197150
rect 123860 197149 126015 197183
rect 123649 197141 126015 197149
rect 125242 197140 126015 197141
rect 123468 197073 123474 197103
rect 123538 197073 123546 197103
rect 123468 197064 123546 197073
rect 123576 197103 123654 197113
rect 123576 197073 123583 197103
rect 123647 197073 123654 197103
rect 123576 196916 123654 197073
rect 123575 196896 123654 196916
rect 123878 197103 123966 197114
rect 123878 197073 123884 197103
rect 123959 197098 123966 197103
rect 123959 197073 123971 197098
rect 123575 196839 123653 196896
rect 123878 196853 123971 197073
rect 123373 196771 123653 196839
rect 123373 196763 123652 196771
rect 122708 196762 123652 196763
rect 121480 196728 123652 196762
rect 121480 196321 123449 196728
rect 123574 196725 123652 196728
rect 121480 196320 122724 196321
rect 101246 193840 101691 193843
rect 121480 195250 121960 196320
rect 122245 196319 122724 196320
rect 101246 193330 101698 193840
rect 121480 193650 121985 195250
rect 123756 193846 124191 196853
rect 125510 195755 126015 197140
rect 145968 197307 146045 197353
rect 145968 197103 146046 197307
rect 148010 197203 148515 197368
rect 146149 197183 148515 197203
rect 146149 197150 146157 197183
rect 146149 197148 146178 197150
rect 146552 197148 148515 197183
rect 146149 197141 148515 197148
rect 145968 197073 145974 197103
rect 146038 197073 146046 197103
rect 145968 197064 146046 197073
rect 146076 197103 146154 197113
rect 146076 197073 146083 197103
rect 146147 197073 146154 197103
rect 146578 197103 146666 197114
rect 146578 197081 146584 197103
rect 146076 196916 146154 197073
rect 146075 196896 146154 196916
rect 146577 197073 146584 197081
rect 146659 197081 146666 197103
rect 146659 197073 146667 197081
rect 146075 196839 146153 196896
rect 146577 196853 146667 197073
rect 145873 196771 146153 196839
rect 145873 196763 146152 196771
rect 145208 196762 146152 196763
rect 143980 196728 146152 196762
rect 143980 196321 145949 196728
rect 146074 196725 146152 196728
rect 143980 196319 145224 196321
rect 143980 196318 144920 196319
rect 143980 195250 144484 196318
rect 123738 193830 124200 193846
rect 123725 192595 124495 193830
rect 143980 193650 144485 195250
rect 146256 193693 146691 196853
rect 148010 195755 148515 197141
rect 146256 193650 146709 193693
rect 146257 193245 146709 193650
rect 55659 174826 56097 174866
rect 55659 174406 56212 174826
rect 55764 174366 56212 174406
rect 55958 174307 56035 174366
rect 55958 174103 56036 174307
rect 58010 174204 58515 174368
rect 78301 174364 78749 174824
rect 57750 174203 58515 174204
rect 56139 174183 58515 174203
rect 56139 174150 56147 174183
rect 56191 174150 58515 174183
rect 56139 174141 58515 174150
rect 55958 174064 55964 174103
rect 56028 174064 56036 174103
rect 55958 174055 56036 174064
rect 56066 174103 56144 174113
rect 56066 174064 56073 174103
rect 56137 174064 56144 174103
rect 56066 173916 56144 174064
rect 56065 173896 56144 173916
rect 56203 174103 56291 174114
rect 56203 174064 56209 174103
rect 56284 174064 56291 174103
rect 56203 174052 56291 174064
rect 56065 173839 56143 173896
rect 55873 173771 56143 173839
rect 56203 173853 56281 174052
rect 56203 173802 56691 173853
rect 55873 173763 56142 173771
rect 55208 173762 56142 173763
rect 53983 173755 54481 173761
rect 54745 173755 56142 173762
rect 53983 173728 56142 173755
rect 56204 173733 56691 173802
rect 53983 173327 55939 173728
rect 56064 173725 56142 173728
rect 56225 173626 56691 173733
rect 53983 172250 54481 173327
rect 54745 173321 55939 173327
rect 54745 173319 55224 173321
rect 53980 170650 54485 172250
rect 56256 170810 56691 173626
rect 58010 172755 58515 174141
rect 78468 174307 78545 174364
rect 78468 174103 78546 174307
rect 80510 174203 81015 174368
rect 100761 174360 101209 174820
rect 78649 174183 81015 174203
rect 78649 174150 78657 174183
rect 78691 174150 81015 174183
rect 78649 174141 81015 174150
rect 78468 174064 78474 174103
rect 78538 174064 78546 174103
rect 78468 174055 78546 174064
rect 78576 174103 78654 174113
rect 78576 174064 78583 174103
rect 78647 174064 78654 174103
rect 78576 173916 78654 174064
rect 78575 173896 78654 173916
rect 78728 174103 78816 174114
rect 78728 174064 78734 174103
rect 78809 174064 78816 174103
rect 78728 174052 78816 174064
rect 78575 173839 78653 173896
rect 78373 173771 78653 173839
rect 78728 173853 78806 174052
rect 78728 173802 79191 173853
rect 76480 173761 76989 173764
rect 78373 173763 78652 173771
rect 77708 173762 78652 173763
rect 77245 173761 78652 173762
rect 76480 173728 78652 173761
rect 78729 173733 79191 173802
rect 76480 173321 78449 173728
rect 78574 173725 78652 173728
rect 76480 173320 77724 173321
rect 76480 172242 76989 173320
rect 77245 173319 77724 173320
rect 56245 170767 56845 170810
rect 56240 170661 56845 170767
rect 56227 170201 56845 170661
rect 76480 170650 76985 172242
rect 78756 170895 79191 173733
rect 80510 172755 81015 174141
rect 100968 174307 101045 174360
rect 100968 174103 101046 174307
rect 103010 174203 103515 174368
rect 123281 174363 123729 174823
rect 101149 174183 103515 174203
rect 101149 174150 101157 174183
rect 101191 174150 103515 174183
rect 101149 174141 103515 174150
rect 100968 174064 100974 174103
rect 101038 174064 101046 174103
rect 100968 174055 101046 174064
rect 101076 174103 101154 174113
rect 101076 174064 101083 174103
rect 101147 174064 101154 174103
rect 101076 173916 101154 174064
rect 101278 174103 101366 174114
rect 101278 174064 101284 174103
rect 101359 174064 101366 174103
rect 101278 174052 101366 174064
rect 101278 174031 101356 174052
rect 101075 173896 101154 173916
rect 101075 173839 101153 173896
rect 101277 173853 101357 174031
rect 100873 173771 101153 173839
rect 100873 173763 101152 173771
rect 100208 173762 101152 173763
rect 99745 173760 101152 173762
rect 99230 173750 101152 173760
rect 98977 173728 101152 173750
rect 101273 173732 101691 173853
rect 98977 173321 100949 173728
rect 101074 173725 101152 173728
rect 98977 172250 99481 173321
rect 99745 173319 100224 173321
rect 98977 172223 99485 172250
rect 78740 170715 79191 170895
rect 56245 169880 56845 170201
rect 78720 169785 79320 170715
rect 98980 170650 99485 172223
rect 101256 170843 101691 173732
rect 103010 172755 103515 174141
rect 123468 174307 123545 174363
rect 123468 174103 123546 174307
rect 125510 174203 126015 174368
rect 145762 174360 146210 174820
rect 123649 174183 126015 174203
rect 123649 174150 123657 174183
rect 123649 174149 123691 174150
rect 123860 174149 126015 174183
rect 123649 174141 126015 174149
rect 125242 174140 126015 174141
rect 123468 174064 123474 174103
rect 123538 174064 123546 174103
rect 123468 174055 123546 174064
rect 123576 174103 123654 174113
rect 123576 174064 123583 174103
rect 123647 174064 123654 174103
rect 123576 173916 123654 174064
rect 123575 173896 123654 173916
rect 123878 174103 123966 174114
rect 123878 174064 123884 174103
rect 123959 174098 123966 174103
rect 123959 174064 123971 174098
rect 123575 173839 123653 173896
rect 123878 173853 123971 174064
rect 123373 173771 123653 173839
rect 123373 173763 123652 173771
rect 122708 173762 123652 173763
rect 121480 173728 123652 173762
rect 121480 173321 123449 173728
rect 123574 173725 123652 173728
rect 121480 173320 122724 173321
rect 101246 170842 101691 170843
rect 101232 170680 101691 170842
rect 121480 172250 121960 173320
rect 122245 173319 122724 173320
rect 101150 169750 101750 170680
rect 121480 170650 121985 172250
rect 123756 170931 124191 173853
rect 125510 172755 126015 174140
rect 145968 174307 146045 174360
rect 145968 174103 146046 174307
rect 148010 174203 148515 174368
rect 146149 174183 148515 174203
rect 146149 174150 146157 174183
rect 146149 174148 146178 174150
rect 146552 174148 148515 174183
rect 146149 174141 148515 174148
rect 145968 174064 145974 174103
rect 146038 174064 146046 174103
rect 145968 174055 146046 174064
rect 146076 174103 146154 174113
rect 146076 174064 146083 174103
rect 146147 174064 146154 174103
rect 146578 174103 146666 174114
rect 146578 174081 146584 174103
rect 146076 173916 146154 174064
rect 146075 173896 146154 173916
rect 146577 174064 146584 174081
rect 146659 174081 146666 174103
rect 146659 174064 146667 174081
rect 146075 173839 146153 173896
rect 146577 173853 146667 174064
rect 145873 173771 146153 173839
rect 145873 173763 146152 173771
rect 145208 173762 146152 173763
rect 143980 173728 146152 173762
rect 143980 173321 145949 173728
rect 146074 173725 146152 173728
rect 143980 173319 145224 173321
rect 143980 173318 144920 173319
rect 143980 172250 144484 173318
rect 123745 170846 124193 170931
rect 123738 170730 124200 170846
rect 123730 169800 124330 170730
rect 143980 170650 144485 172250
rect 146256 170860 146691 173853
rect 148010 172755 148515 174141
rect 146256 170837 147130 170860
rect 146232 170745 147130 170837
rect 146085 169930 147130 170745
rect 146085 169815 146685 169930
rect 78258 152246 78725 152252
rect 55906 151368 56246 151572
rect 78258 151371 78726 152246
rect 100900 151982 101231 152005
rect 55958 151307 56035 151368
rect 55958 151103 56036 151307
rect 58010 151204 58515 151368
rect 78259 151365 78726 151371
rect 100894 151373 101231 151982
rect 57750 151203 58515 151204
rect 56139 151183 58515 151203
rect 56139 151150 56147 151183
rect 56191 151150 58515 151183
rect 56139 151141 58515 151150
rect 55958 151044 55964 151103
rect 56028 151044 56036 151103
rect 55958 151035 56036 151044
rect 56066 151103 56144 151113
rect 56066 151044 56073 151103
rect 56137 151044 56144 151103
rect 56066 150916 56144 151044
rect 56065 150896 56144 150916
rect 56203 151103 56291 151114
rect 56203 151044 56209 151103
rect 56284 151044 56291 151103
rect 56203 151032 56291 151044
rect 56065 150839 56143 150896
rect 55873 150771 56143 150839
rect 56203 150853 56281 151032
rect 56203 150802 56691 150853
rect 55873 150763 56142 150771
rect 55208 150762 56142 150763
rect 53983 150755 54481 150761
rect 54745 150755 56142 150762
rect 53983 150728 56142 150755
rect 56204 150733 56691 150802
rect 53983 150327 55939 150728
rect 56064 150725 56142 150728
rect 56225 150626 56691 150733
rect 53983 149250 54481 150327
rect 54745 150321 55939 150327
rect 54745 150319 55224 150321
rect 53980 147650 54485 149250
rect 56256 148022 56691 150626
rect 58010 149755 58515 151141
rect 78468 151307 78545 151365
rect 78468 151103 78546 151307
rect 80510 151203 81015 151368
rect 100894 151350 101225 151373
rect 78649 151183 81015 151203
rect 78649 151150 78657 151183
rect 78691 151150 81015 151183
rect 78649 151141 81015 151150
rect 78468 151044 78474 151103
rect 78538 151044 78546 151103
rect 78468 151035 78546 151044
rect 78576 151103 78654 151113
rect 78576 151044 78583 151103
rect 78647 151044 78654 151103
rect 78576 150916 78654 151044
rect 78575 150896 78654 150916
rect 78728 151103 78816 151114
rect 78728 151044 78734 151103
rect 78809 151044 78816 151103
rect 78728 151032 78816 151044
rect 78575 150839 78653 150896
rect 78373 150771 78653 150839
rect 78728 150853 78806 151032
rect 78728 150802 79191 150853
rect 76480 150761 76989 150764
rect 78373 150763 78652 150771
rect 77708 150762 78652 150763
rect 77245 150761 78652 150762
rect 76480 150728 78652 150761
rect 78729 150733 79191 150802
rect 76480 150321 78449 150728
rect 78574 150725 78652 150728
rect 76480 150320 77724 150321
rect 76480 149242 76989 150320
rect 77245 150319 77724 150320
rect 56229 147767 56693 148022
rect 56229 147650 56696 147767
rect 76480 147650 76985 149242
rect 78756 148061 79191 150733
rect 80510 149755 81015 151141
rect 100968 151307 101045 151350
rect 100968 151103 101046 151307
rect 103010 151203 103515 151368
rect 123165 151352 123627 152033
rect 145856 151368 146232 151719
rect 101149 151183 103515 151203
rect 101149 151150 101157 151183
rect 101191 151150 103515 151183
rect 101149 151141 103515 151150
rect 100968 151044 100974 151103
rect 101038 151044 101046 151103
rect 100968 151035 101046 151044
rect 101076 151103 101154 151113
rect 101076 151044 101083 151103
rect 101147 151044 101154 151103
rect 101076 150916 101154 151044
rect 101278 151103 101366 151114
rect 101278 151044 101284 151103
rect 101359 151044 101366 151103
rect 101278 151032 101366 151044
rect 101278 151031 101364 151032
rect 101075 150896 101154 150916
rect 101277 151015 101364 151031
rect 101075 150839 101153 150896
rect 101277 150853 101357 151015
rect 100873 150771 101153 150839
rect 100873 150763 101152 150771
rect 100208 150762 101152 150763
rect 99745 150760 101152 150762
rect 99230 150750 101152 150760
rect 98977 150728 101152 150750
rect 101273 150732 101691 150853
rect 98977 150321 100949 150728
rect 101074 150725 101152 150728
rect 98977 149250 99481 150321
rect 99745 150319 100224 150321
rect 98977 149223 99485 149250
rect 78746 147815 79213 148061
rect 78744 147650 79213 147815
rect 98980 147650 99485 149223
rect 101256 147966 101691 150732
rect 103010 149755 103515 151141
rect 123468 151307 123545 151352
rect 123468 151103 123546 151307
rect 125510 151203 126015 151368
rect 123649 151183 126015 151203
rect 123649 151150 123657 151183
rect 123649 151149 123691 151150
rect 123860 151149 126015 151183
rect 123649 151141 126015 151149
rect 125242 151140 126015 151141
rect 123468 151044 123474 151103
rect 123538 151044 123546 151103
rect 123468 151035 123546 151044
rect 123576 151103 123654 151113
rect 123576 151044 123583 151103
rect 123647 151044 123654 151103
rect 123576 150916 123654 151044
rect 123575 150896 123654 150916
rect 123878 151103 123966 151114
rect 123878 151044 123884 151103
rect 123959 151098 123966 151103
rect 123959 151044 123971 151098
rect 123575 150839 123653 150896
rect 123878 150853 123971 151044
rect 123373 150771 123653 150839
rect 123373 150763 123652 150771
rect 122708 150762 123652 150763
rect 121480 150728 123652 150762
rect 121480 150321 123449 150728
rect 123574 150725 123652 150728
rect 121480 150320 122724 150321
rect 121480 149250 121960 150320
rect 122245 150319 122724 150320
rect 56229 147223 56693 147650
rect 78746 147180 79213 147650
rect 101223 146997 101724 147966
rect 121480 147650 121985 149250
rect 123756 147946 124191 150853
rect 125510 149755 126015 151140
rect 145968 151307 146045 151368
rect 145968 151103 146046 151307
rect 148010 151203 148515 151368
rect 146149 151183 148515 151203
rect 146149 151150 146157 151183
rect 146149 151148 146178 151150
rect 146552 151148 148515 151183
rect 146149 151141 148515 151148
rect 145968 151044 145974 151103
rect 146038 151044 146046 151103
rect 145968 151035 146046 151044
rect 146076 151103 146154 151113
rect 146076 151044 146083 151103
rect 146147 151044 146154 151103
rect 146578 151103 146666 151114
rect 146578 151081 146584 151103
rect 146076 150916 146154 151044
rect 146075 150896 146154 150916
rect 146577 151044 146584 151081
rect 146659 151081 146666 151103
rect 146659 151044 146667 151081
rect 146075 150839 146153 150896
rect 146577 150853 146667 151044
rect 145873 150771 146153 150839
rect 145873 150763 146152 150771
rect 145208 150762 146152 150763
rect 143980 150728 146152 150762
rect 143980 150321 145949 150728
rect 146074 150725 146152 150728
rect 143980 150319 145224 150321
rect 143980 150318 144920 150319
rect 143980 149250 144484 150318
rect 123756 147846 124220 147946
rect 123738 147650 124220 147846
rect 143980 147650 144485 149250
rect 146256 148078 146691 150853
rect 148010 149755 148515 151141
rect 123758 147295 124220 147650
rect 146204 146975 146691 148078
rect 55817 128367 56265 128939
rect 55958 128307 56035 128367
rect 55958 128103 56036 128307
rect 58010 128204 58515 128368
rect 78291 128351 78739 128923
rect 57750 128203 58515 128204
rect 56139 128183 58515 128203
rect 56139 128150 56147 128183
rect 56191 128150 58515 128183
rect 56139 128141 58515 128150
rect 55958 128028 55964 128103
rect 56028 128028 56036 128103
rect 55958 128019 56036 128028
rect 56066 128103 56144 128113
rect 56066 128028 56073 128103
rect 56137 128028 56144 128103
rect 56066 127916 56144 128028
rect 56065 127896 56144 127916
rect 56203 128103 56291 128114
rect 56203 128028 56209 128103
rect 56284 128028 56291 128103
rect 56203 128016 56291 128028
rect 56065 127839 56143 127896
rect 55873 127771 56143 127839
rect 56203 127853 56281 128016
rect 56203 127802 56691 127853
rect 55873 127763 56142 127771
rect 55208 127762 56142 127763
rect 53983 127755 54481 127761
rect 54745 127755 56142 127762
rect 53983 127728 56142 127755
rect 56204 127733 56691 127802
rect 53983 127327 55939 127728
rect 56064 127725 56142 127728
rect 56225 127626 56691 127733
rect 53983 126250 54481 127327
rect 54745 127321 55939 127327
rect 54745 127319 55224 127321
rect 53980 124650 54485 126250
rect 56256 125025 56691 127626
rect 58010 126755 58515 128141
rect 78468 128307 78545 128351
rect 78468 128103 78546 128307
rect 80510 128203 81015 128368
rect 100767 128361 101215 128946
rect 78649 128183 81015 128203
rect 78649 128150 78657 128183
rect 78691 128150 81015 128183
rect 78649 128141 81015 128150
rect 78468 128028 78474 128103
rect 78538 128028 78546 128103
rect 78468 128019 78546 128028
rect 78576 128103 78654 128113
rect 78576 128028 78583 128103
rect 78647 128028 78654 128103
rect 78576 127916 78654 128028
rect 78575 127896 78654 127916
rect 78728 128103 78816 128114
rect 78728 128028 78734 128103
rect 78809 128028 78816 128103
rect 78728 128016 78816 128028
rect 78575 127839 78653 127896
rect 78373 127771 78653 127839
rect 78728 127853 78806 128016
rect 78728 127802 79191 127853
rect 76480 127761 76989 127764
rect 78373 127763 78652 127771
rect 77708 127762 78652 127763
rect 77245 127761 78652 127762
rect 76480 127728 78652 127761
rect 78729 127733 79191 127802
rect 76480 127321 78449 127728
rect 78574 127725 78652 127728
rect 76480 127320 77724 127321
rect 76480 126242 76989 127320
rect 77245 127319 77724 127320
rect 56070 124140 56820 125025
rect 76480 124650 76985 126242
rect 78756 124907 79191 127733
rect 80510 126755 81015 128141
rect 100968 128307 101045 128361
rect 100968 128103 101046 128307
rect 103010 128203 103515 128368
rect 123305 128360 123753 128932
rect 101149 128183 103515 128203
rect 101149 128150 101157 128183
rect 101191 128150 103515 128183
rect 101149 128141 103515 128150
rect 100968 128028 100974 128103
rect 101038 128028 101046 128103
rect 100968 128019 101046 128028
rect 101076 128103 101154 128113
rect 101076 128028 101083 128103
rect 101147 128028 101154 128103
rect 101278 128103 101366 128114
rect 101278 128031 101284 128103
rect 101076 127916 101154 128028
rect 101075 127896 101154 127916
rect 101277 128028 101284 128031
rect 101359 128028 101366 128103
rect 101277 128016 101366 128028
rect 101075 127839 101153 127896
rect 101277 127853 101357 128016
rect 100873 127771 101153 127839
rect 100873 127763 101152 127771
rect 100208 127762 101152 127763
rect 99745 127760 101152 127762
rect 99230 127750 101152 127760
rect 98977 127728 101152 127750
rect 101273 127732 101691 127853
rect 98977 127321 100949 127728
rect 101074 127725 101152 127728
rect 98977 126250 99481 127321
rect 99745 127319 100224 127321
rect 98977 126223 99485 126250
rect 78751 124815 79199 124907
rect 78744 124650 79199 124815
rect 98980 124650 99485 126223
rect 101256 124843 101691 127732
rect 103010 126755 103515 128141
rect 123468 128307 123545 128360
rect 123468 128103 123546 128307
rect 125510 128203 126015 128368
rect 145780 128345 146228 128917
rect 123649 128183 126015 128203
rect 123649 128150 123657 128183
rect 123649 128149 123691 128150
rect 123860 128149 126015 128183
rect 123649 128141 126015 128149
rect 125242 128140 126015 128141
rect 123468 128028 123474 128103
rect 123538 128028 123546 128103
rect 123468 128019 123546 128028
rect 123576 128103 123654 128113
rect 123576 128028 123583 128103
rect 123647 128028 123654 128103
rect 123576 127916 123654 128028
rect 123575 127896 123654 127916
rect 123878 128103 123966 128114
rect 123878 128028 123884 128103
rect 123959 128098 123966 128103
rect 123959 128028 123971 128098
rect 123575 127839 123653 127896
rect 123878 127853 123971 128028
rect 123373 127771 123653 127839
rect 123373 127763 123652 127771
rect 122708 127762 123652 127763
rect 121480 127728 123652 127762
rect 121480 127321 123449 127728
rect 123574 127725 123652 127728
rect 121480 127320 122724 127321
rect 101246 124781 101691 124843
rect 121480 126250 121960 127320
rect 122245 127319 122724 127320
rect 101246 124650 101699 124781
rect 121480 124650 121985 126250
rect 123756 124970 124191 127853
rect 125510 126755 126015 128140
rect 145968 128307 146045 128345
rect 145968 128103 146046 128307
rect 148010 128203 148515 128368
rect 146149 128183 148515 128203
rect 146149 128150 146157 128183
rect 146149 128148 146178 128150
rect 146552 128148 148515 128183
rect 146149 128141 148515 128148
rect 145968 128028 145974 128103
rect 146038 128028 146046 128103
rect 145968 128019 146046 128028
rect 146076 128103 146154 128113
rect 146076 128028 146083 128103
rect 146147 128028 146154 128103
rect 146578 128103 146666 128114
rect 146578 128081 146584 128103
rect 146076 127916 146154 128028
rect 146075 127896 146154 127916
rect 146577 128028 146584 128081
rect 146659 128081 146666 128103
rect 146659 128028 146667 128081
rect 146075 127839 146153 127896
rect 146577 127853 146667 128028
rect 145873 127771 146153 127839
rect 145873 127763 146152 127771
rect 145208 127762 146152 127763
rect 143980 127728 146152 127762
rect 143980 127321 145949 127728
rect 146074 127725 146152 127728
rect 143980 127319 145224 127321
rect 143980 127318 144920 127319
rect 143980 126250 144484 127318
rect 123756 124846 124205 124970
rect 123738 124775 124205 124846
rect 78751 124335 79199 124650
rect 101251 124209 101699 124650
rect 123695 123845 124295 124775
rect 143980 124650 144485 126250
rect 146256 124728 146691 127853
rect 148010 126755 148515 128141
rect 146255 124156 146703 124728
rect 145717 105995 146147 106013
rect 55800 105352 56230 105992
rect 55958 105307 56035 105352
rect 55958 105103 56036 105307
rect 58010 105204 58515 105368
rect 78289 105346 78719 105986
rect 57750 105203 58515 105204
rect 56139 105183 58515 105203
rect 56139 105150 56147 105183
rect 56191 105150 58515 105183
rect 56139 105141 58515 105150
rect 55958 104963 55964 105103
rect 56028 104963 56036 105103
rect 55958 104954 56036 104963
rect 56066 105103 56144 105113
rect 56066 104963 56073 105103
rect 56137 104963 56144 105103
rect 56066 104916 56144 104963
rect 56065 104896 56144 104916
rect 56203 105103 56291 105114
rect 56203 104963 56209 105103
rect 56284 104963 56291 105103
rect 56203 104951 56291 104963
rect 56065 104839 56143 104896
rect 55873 104771 56143 104839
rect 56203 104853 56281 104951
rect 56203 104802 56691 104853
rect 55873 104763 56142 104771
rect 55208 104762 56142 104763
rect 53983 104755 54481 104761
rect 54745 104755 56142 104762
rect 53983 104728 56142 104755
rect 56204 104733 56691 104802
rect 53983 104327 55939 104728
rect 56064 104725 56142 104728
rect 56225 104626 56691 104733
rect 53983 103250 54481 104327
rect 54745 104321 55939 104327
rect 54745 104319 55224 104321
rect 53980 101650 54485 103250
rect 56256 101957 56691 104626
rect 58010 103755 58515 105141
rect 78468 105307 78545 105346
rect 78468 105103 78546 105307
rect 80510 105203 81015 105368
rect 100759 105355 101189 105995
rect 78649 105183 81015 105203
rect 78649 105150 78657 105183
rect 78691 105150 81015 105183
rect 78649 105141 81015 105150
rect 78468 104963 78474 105103
rect 78538 104963 78546 105103
rect 78468 104954 78546 104963
rect 78576 105103 78654 105113
rect 78576 104963 78583 105103
rect 78647 104963 78654 105103
rect 78576 104916 78654 104963
rect 78575 104896 78654 104916
rect 78728 105103 78816 105114
rect 78728 104963 78734 105103
rect 78809 104963 78816 105103
rect 78728 104951 78816 104963
rect 78575 104839 78653 104896
rect 78373 104771 78653 104839
rect 78728 104853 78806 104951
rect 78728 104802 79191 104853
rect 76480 104761 76989 104764
rect 78373 104763 78652 104771
rect 77708 104762 78652 104763
rect 77245 104761 78652 104762
rect 76480 104728 78652 104761
rect 78729 104733 79191 104802
rect 76480 104321 78449 104728
rect 78574 104725 78652 104728
rect 76480 104320 77724 104321
rect 76480 103242 76989 104320
rect 77245 104319 77724 104320
rect 56256 101767 56714 101957
rect 56240 101650 56714 101767
rect 76480 101650 76985 103242
rect 78756 101859 79191 104733
rect 80510 103755 81015 105141
rect 100968 105307 101045 105355
rect 100968 105103 101046 105307
rect 103010 105203 103515 105368
rect 123238 105346 123668 105986
rect 145708 105373 146147 105995
rect 101149 105183 103515 105203
rect 101149 105150 101157 105183
rect 101191 105150 103515 105183
rect 101149 105141 103515 105150
rect 100968 104963 100974 105103
rect 101038 104963 101046 105103
rect 100968 104954 101046 104963
rect 101076 105103 101154 105113
rect 101076 104963 101083 105103
rect 101147 104963 101154 105103
rect 101278 105103 101366 105114
rect 101278 105031 101284 105103
rect 101076 104916 101154 104963
rect 101075 104896 101154 104916
rect 101277 104963 101284 105031
rect 101359 104963 101366 105103
rect 101277 104951 101366 104963
rect 101075 104839 101153 104896
rect 101277 104853 101357 104951
rect 100873 104771 101153 104839
rect 100873 104763 101152 104771
rect 100208 104762 101152 104763
rect 99745 104760 101152 104762
rect 99230 104750 101152 104760
rect 98977 104728 101152 104750
rect 101273 104732 101691 104853
rect 98977 104321 100949 104728
rect 101074 104725 101152 104728
rect 98977 103250 99481 104321
rect 99745 104319 100224 104321
rect 98977 103223 99485 103250
rect 78756 101815 79196 101859
rect 78744 101650 79196 101815
rect 98980 101650 99485 103223
rect 101256 101843 101691 104732
rect 103010 103755 103515 105141
rect 123468 105307 123545 105346
rect 123468 105103 123546 105307
rect 125510 105203 126015 105368
rect 145708 105355 146138 105373
rect 123649 105183 126015 105203
rect 123649 105150 123657 105183
rect 123649 105149 123691 105150
rect 123860 105149 126015 105183
rect 123649 105141 126015 105149
rect 125242 105140 126015 105141
rect 123468 104963 123474 105103
rect 123538 104963 123546 105103
rect 123468 104954 123546 104963
rect 123576 105103 123654 105113
rect 123576 104963 123583 105103
rect 123647 104963 123654 105103
rect 123576 104916 123654 104963
rect 123575 104896 123654 104916
rect 123878 105103 123966 105114
rect 123878 104963 123884 105103
rect 123959 105098 123966 105103
rect 123959 104963 123971 105098
rect 123575 104839 123653 104896
rect 123878 104853 123971 104963
rect 123373 104771 123653 104839
rect 123373 104763 123652 104771
rect 122708 104762 123652 104763
rect 121480 104728 123652 104762
rect 121480 104321 123449 104728
rect 123574 104725 123652 104728
rect 121480 104320 122724 104321
rect 101246 101841 101691 101843
rect 101245 101650 101691 101841
rect 121480 103250 121960 104320
rect 122245 104319 122724 104320
rect 121480 101650 121985 103250
rect 123756 101846 124191 104853
rect 125510 103755 126015 105140
rect 145968 105307 146045 105355
rect 145968 105103 146046 105307
rect 148010 105203 148515 105368
rect 146149 105183 148515 105203
rect 146149 105150 146157 105183
rect 146149 105148 146178 105150
rect 146552 105148 148515 105183
rect 146149 105141 148515 105148
rect 145968 104963 145974 105103
rect 146038 104963 146046 105103
rect 145968 104954 146046 104963
rect 146076 105103 146154 105113
rect 146076 104963 146083 105103
rect 146147 104963 146154 105103
rect 146578 105103 146666 105114
rect 146578 105081 146584 105103
rect 146076 104916 146154 104963
rect 146075 104896 146154 104916
rect 146577 104963 146584 105081
rect 146659 105081 146666 105103
rect 146659 104963 146667 105081
rect 146075 104839 146153 104896
rect 146577 104853 146667 104963
rect 145873 104771 146153 104839
rect 145873 104763 146152 104771
rect 145208 104762 146152 104763
rect 143980 104728 146152 104762
rect 143980 104321 145949 104728
rect 146074 104725 146152 104728
rect 143980 104319 145224 104321
rect 143980 104318 144920 104319
rect 143980 103250 144484 104318
rect 123738 101650 124200 101846
rect 143980 101650 144485 103250
rect 146256 101706 146691 104853
rect 148010 103755 148515 105141
rect 146221 101650 146691 101706
rect 56266 101317 56714 101650
rect 56266 101313 56696 101317
rect 78766 101219 79196 101650
rect 101245 101201 101675 101650
rect 123742 101201 124172 101650
rect 146221 101066 146651 101650
rect 55807 82344 56247 82899
rect 55958 82307 56035 82344
rect 55958 82103 56036 82307
rect 58010 82204 58515 82368
rect 78184 82344 78624 82899
rect 57750 82203 58515 82204
rect 56139 82183 58515 82203
rect 56139 82150 56147 82183
rect 56191 82150 58515 82183
rect 56139 82141 58515 82150
rect 55958 81839 55964 82103
rect 55873 81828 55964 81839
rect 56028 81839 56036 82103
rect 56066 82103 56144 82113
rect 56066 81916 56073 82103
rect 56065 81839 56073 81916
rect 56028 81828 56073 81839
rect 56137 81828 56144 82103
rect 55873 81816 56144 81828
rect 56203 82103 56291 82114
rect 56203 81828 56209 82103
rect 56284 81853 56291 82103
rect 56284 81828 56691 81853
rect 55873 81771 56143 81816
rect 56203 81802 56691 81828
rect 55873 81763 56142 81771
rect 55208 81762 56142 81763
rect 53983 81755 54481 81761
rect 54745 81755 56142 81762
rect 53983 81728 56142 81755
rect 56204 81733 56691 81802
rect 53983 81327 55939 81728
rect 56064 81725 56142 81728
rect 56225 81626 56691 81733
rect 53983 80250 54481 81327
rect 54745 81321 55939 81327
rect 54745 81319 55224 81321
rect 53980 78650 54485 80250
rect 56256 78810 56691 81626
rect 58010 80755 58515 82141
rect 78468 82307 78545 82344
rect 78468 82103 78546 82307
rect 80510 82203 81015 82368
rect 100755 82362 101195 82917
rect 78649 82183 81015 82203
rect 78649 82150 78657 82183
rect 78691 82150 81015 82183
rect 78649 82141 81015 82150
rect 78468 81839 78474 82103
rect 78373 81828 78474 81839
rect 78538 81839 78546 82103
rect 78576 82103 78654 82113
rect 78576 81916 78583 82103
rect 78575 81839 78583 81916
rect 78538 81828 78583 81839
rect 78647 81828 78654 82103
rect 78373 81816 78654 81828
rect 78728 82103 78816 82114
rect 78728 81828 78734 82103
rect 78809 81853 78816 82103
rect 78809 81828 79191 81853
rect 78373 81771 78653 81816
rect 78728 81802 79191 81828
rect 76480 81761 76989 81764
rect 78373 81763 78652 81771
rect 77708 81762 78652 81763
rect 77245 81761 78652 81762
rect 76480 81728 78652 81761
rect 78729 81733 79191 81802
rect 76480 81321 78449 81728
rect 78574 81725 78652 81728
rect 76480 81320 77724 81321
rect 56213 78767 56691 78810
rect 76480 80242 76989 81320
rect 77245 81319 77724 81320
rect 56213 78650 56696 78767
rect 76480 78650 76985 80242
rect 78756 78871 79191 81733
rect 80510 80755 81015 82141
rect 100968 82307 101045 82362
rect 100968 82103 101046 82307
rect 103010 82203 103515 82368
rect 123273 82353 123713 82908
rect 101149 82183 103515 82203
rect 101149 82150 101157 82183
rect 101191 82150 103515 82183
rect 101149 82141 103515 82150
rect 100968 81839 100974 82103
rect 100873 81828 100974 81839
rect 101038 81839 101046 82103
rect 101076 82103 101154 82113
rect 101076 81916 101083 82103
rect 101075 81839 101083 81916
rect 101038 81828 101083 81839
rect 101147 81828 101154 82103
rect 101278 82103 101366 82114
rect 101278 82031 101284 82103
rect 101277 81853 101284 82031
rect 100873 81816 101154 81828
rect 101273 81828 101284 81853
rect 101359 81853 101366 82103
rect 101359 81828 101691 81853
rect 100873 81771 101153 81816
rect 100873 81763 101152 81771
rect 100208 81762 101152 81763
rect 99745 81760 101152 81762
rect 99230 81750 101152 81760
rect 98977 81728 101152 81750
rect 101273 81732 101691 81828
rect 98977 81321 100949 81728
rect 101074 81725 101152 81728
rect 98977 80250 99481 81321
rect 99745 81319 100224 81321
rect 98977 80223 99485 80250
rect 78740 78650 79191 78871
rect 98980 78650 99485 80223
rect 101256 78843 101691 81732
rect 103010 80755 103515 82141
rect 123468 82307 123545 82353
rect 123468 82103 123546 82307
rect 125510 82203 126015 82368
rect 145659 82344 146099 82899
rect 123649 82183 126015 82203
rect 123649 82150 123657 82183
rect 123649 82149 123691 82150
rect 123860 82149 126015 82183
rect 123649 82141 126015 82149
rect 125242 82140 126015 82141
rect 123468 81839 123474 82103
rect 123373 81828 123474 81839
rect 123538 81839 123546 82103
rect 123576 82103 123654 82113
rect 123576 81916 123583 82103
rect 123575 81839 123583 81916
rect 123538 81828 123583 81839
rect 123647 81828 123654 82103
rect 123878 82103 123966 82114
rect 123878 81853 123884 82103
rect 123373 81816 123654 81828
rect 123756 81828 123884 81853
rect 123959 82098 123966 82103
rect 123959 81853 123971 82098
rect 123959 81828 124191 81853
rect 123373 81771 123653 81816
rect 123373 81763 123652 81771
rect 122708 81762 123652 81763
rect 121480 81728 123652 81762
rect 121480 81321 123449 81728
rect 123574 81725 123652 81728
rect 121480 81320 122724 81321
rect 101246 78775 101691 78843
rect 101231 78650 101691 78775
rect 121480 80250 121960 81320
rect 122245 81319 122724 81320
rect 121480 78650 121985 80250
rect 123756 78846 124191 81828
rect 125510 80755 126015 82140
rect 145968 82307 146045 82344
rect 145968 82103 146046 82307
rect 148010 82203 148515 82368
rect 146149 82183 148515 82203
rect 146149 82150 146157 82183
rect 146149 82148 146178 82150
rect 146552 82148 148515 82183
rect 146149 82141 148515 82148
rect 145968 81839 145974 82103
rect 145873 81828 145974 81839
rect 146038 81839 146046 82103
rect 146076 82103 146154 82113
rect 146076 81916 146083 82103
rect 146075 81839 146083 81916
rect 146038 81828 146083 81839
rect 146147 81828 146154 82103
rect 146578 82103 146666 82114
rect 146578 82081 146584 82103
rect 146577 81853 146584 82081
rect 145873 81816 146154 81828
rect 146256 81828 146584 81853
rect 146659 82081 146666 82103
rect 146659 81853 146667 82081
rect 146659 81828 146691 81853
rect 145873 81771 146153 81816
rect 145873 81763 146152 81771
rect 145208 81762 146152 81763
rect 143980 81728 146152 81762
rect 143980 81321 145949 81728
rect 146074 81725 146152 81728
rect 143980 81319 145224 81321
rect 143980 81318 144920 81319
rect 143980 80250 144484 81318
rect 123738 78819 124200 78846
rect 123738 78650 124216 78819
rect 143980 78650 144485 80250
rect 146256 78827 146691 81828
rect 148010 80755 148515 82141
rect 146250 78650 146691 78827
rect 56213 78255 56653 78650
rect 78740 78316 79180 78650
rect 101231 78220 101671 78650
rect 123776 78264 124216 78650
rect 146250 78272 146690 78650
rect 55667 59365 56218 59608
rect 55958 59307 56035 59365
rect 55958 59103 56036 59307
rect 58010 59204 58515 59368
rect 78358 59359 78746 59616
rect 57750 59203 58515 59204
rect 56139 59183 58515 59203
rect 56139 59150 56147 59183
rect 56191 59150 58515 59183
rect 56139 59141 58515 59150
rect 55208 58762 55657 58763
rect 53983 58755 54481 58761
rect 54745 58755 55657 58762
rect 53983 58560 55657 58755
rect 55958 58628 55964 59103
rect 56028 58628 56036 59103
rect 55958 58619 56036 58628
rect 56066 59103 56144 59113
rect 56066 58628 56073 59103
rect 56137 58628 56144 59103
rect 56066 58560 56144 58628
rect 56203 59103 56291 59114
rect 56203 58628 56209 59103
rect 56284 58997 56291 59103
rect 56284 58853 56568 58997
rect 56284 58628 56691 58853
rect 56203 58616 56691 58628
rect 53983 58327 56149 58560
rect 53983 57250 54481 58327
rect 54745 58321 56149 58327
rect 54745 58319 55224 58321
rect 55608 58317 56149 58321
rect 53980 55650 54485 57250
rect 56256 55840 56691 58616
rect 58010 57755 58515 59141
rect 78468 59307 78545 59359
rect 78468 59103 78546 59307
rect 80510 59203 81015 59368
rect 100865 59352 101246 59639
rect 78649 59183 81015 59203
rect 78649 59150 78657 59183
rect 78691 59150 81015 59183
rect 78649 59141 81015 59150
rect 76480 58761 76989 58764
rect 77708 58762 78121 58763
rect 77245 58761 78121 58762
rect 76480 58557 78121 58761
rect 78468 58628 78474 59103
rect 78538 58628 78546 59103
rect 78576 59103 78654 59113
rect 78576 58916 78583 59103
rect 78575 58725 78583 58916
rect 78468 58619 78546 58628
rect 78576 58628 78583 58725
rect 78647 58628 78654 59103
rect 78576 58557 78654 58628
rect 78728 59103 78816 59114
rect 78728 58628 78734 59103
rect 78809 58992 78816 59103
rect 78809 58853 78980 58992
rect 78809 58628 79191 58853
rect 78728 58616 79191 58628
rect 76480 58321 78654 58557
rect 76480 58320 77724 58321
rect 76480 57242 76989 58320
rect 77245 58319 77724 58320
rect 56225 55830 56825 55840
rect 56160 54910 56825 55830
rect 76480 55650 76985 57242
rect 78756 55815 79191 58616
rect 80510 57755 81015 59141
rect 100968 59307 101045 59352
rect 100968 59103 101046 59307
rect 103010 59203 103515 59368
rect 123331 59353 123714 59685
rect 101149 59183 103515 59203
rect 101149 59150 101157 59183
rect 101191 59150 103515 59183
rect 101149 59141 103515 59150
rect 100208 58762 100539 58763
rect 99745 58760 100539 58762
rect 99230 58750 100539 58760
rect 98977 58561 100539 58750
rect 100968 58628 100974 59103
rect 101038 58628 101046 59103
rect 101076 59103 101154 59113
rect 101076 58916 101083 59103
rect 101075 58725 101083 58916
rect 100968 58619 101046 58628
rect 101076 58628 101083 58725
rect 101147 58628 101154 59103
rect 101278 59103 101366 59114
rect 101278 59031 101284 59103
rect 101277 58853 101284 59031
rect 101273 58732 101284 58853
rect 101076 58561 101154 58628
rect 98977 58509 101154 58561
rect 101256 58628 101284 58732
rect 101359 58853 101366 59103
rect 101359 58628 101691 58853
rect 98977 58321 101153 58509
rect 98977 57250 99481 58321
rect 99745 58319 100224 58321
rect 100509 58318 101153 58321
rect 98977 57223 99485 57250
rect 78744 55800 79191 55815
rect 56160 54900 56760 54910
rect 78670 54870 79270 55800
rect 98980 55650 99485 57223
rect 101256 56073 101691 58628
rect 103010 57755 103515 59141
rect 123468 59307 123545 59353
rect 123468 59103 123546 59307
rect 125510 59203 126015 59368
rect 145772 59361 146246 59789
rect 123649 59183 126015 59203
rect 123649 59150 123657 59183
rect 123649 59149 123691 59150
rect 123860 59149 126015 59183
rect 123649 59141 126015 59149
rect 125242 59140 126015 59141
rect 122708 58762 123196 58763
rect 121480 58561 123196 58762
rect 123468 58628 123474 59103
rect 123538 58628 123546 59103
rect 123576 59103 123654 59113
rect 123576 58916 123583 59103
rect 123575 58725 123583 58916
rect 123468 58619 123546 58628
rect 123576 58628 123583 58725
rect 123647 58628 123654 59103
rect 123878 59103 123966 59114
rect 123878 58853 123884 59103
rect 123576 58561 123654 58628
rect 121480 58478 123654 58561
rect 123877 58628 123884 58853
rect 123959 59098 123966 59103
rect 123959 58853 123971 59098
rect 123959 58628 124191 58853
rect 121480 58321 123651 58478
rect 121480 58320 122724 58321
rect 121480 57250 121960 58320
rect 122245 58319 122724 58320
rect 123039 58316 123651 58321
rect 123877 58115 124191 58628
rect 101244 55855 101696 56073
rect 101244 55298 101880 55855
rect 121480 55650 121985 57250
rect 123756 55912 124191 58115
rect 125510 57755 126015 59140
rect 145968 59307 146045 59361
rect 145968 59103 146046 59307
rect 148010 59203 148515 59368
rect 146149 59183 148515 59203
rect 146149 59150 146157 59183
rect 146149 59148 146178 59150
rect 146552 59148 148515 59183
rect 146149 59141 148515 59148
rect 145208 58762 145562 58763
rect 143980 58541 145562 58762
rect 145968 58628 145974 59103
rect 146038 58628 146046 59103
rect 146076 59103 146154 59113
rect 146076 58916 146083 59103
rect 146075 58725 146083 58916
rect 145968 58619 146046 58628
rect 146076 58628 146083 58725
rect 146147 58628 146154 59103
rect 146578 59103 146666 59114
rect 146578 59081 146584 59103
rect 146076 58541 146154 58628
rect 143980 58525 146154 58541
rect 146577 58628 146584 59081
rect 146659 59081 146666 59103
rect 146659 58853 146667 59081
rect 146659 58628 146691 58853
rect 143980 58324 146151 58525
rect 143980 58321 145562 58324
rect 143980 58319 145224 58321
rect 143980 58318 144920 58319
rect 143980 57250 144484 58318
rect 146577 58044 146691 58628
rect 123581 55421 124385 55912
rect 143980 55650 144485 57250
rect 146256 55844 146691 58044
rect 148010 57755 148515 59141
rect 146242 55695 146716 55844
rect 101280 54925 101880 55298
rect 123685 54790 124285 55421
rect 146230 54765 146830 55695
rect 55837 36363 56211 36787
rect 55958 36307 56035 36363
rect 55958 36103 56036 36307
rect 58010 36204 58515 36368
rect 78194 36354 78691 36837
rect 57750 36203 58515 36204
rect 56139 36183 58515 36203
rect 56139 36150 56147 36183
rect 56191 36150 58515 36183
rect 56139 36141 58515 36150
rect 55958 35428 55964 36103
rect 56028 35428 56036 36103
rect 55958 35419 56036 35428
rect 56066 36103 56144 36113
rect 56066 35428 56073 36103
rect 56137 35428 56144 36103
rect 56066 35416 56144 35428
rect 56203 36103 56291 36114
rect 56203 35428 56209 36103
rect 56284 35865 56291 36103
rect 56284 35428 56618 35865
rect 56203 35416 56618 35428
rect 58010 35416 58515 36141
rect 78468 36307 78545 36354
rect 78468 36103 78546 36307
rect 80510 36203 81015 36368
rect 100777 36361 101214 36702
rect 78649 36183 81015 36203
rect 78649 36150 78657 36183
rect 78691 36150 81015 36183
rect 78649 36141 81015 36150
rect 78468 35428 78474 36103
rect 78538 35428 78546 36103
rect 78576 36103 78654 36113
rect 78576 35554 78583 36103
rect 78468 35419 78546 35428
rect 78575 35428 78583 35554
rect 78647 35428 78654 36103
rect 78575 35416 78654 35428
rect 78728 36103 78816 36114
rect 78728 35428 78734 36103
rect 78809 35757 78816 36103
rect 78809 35428 79001 35757
rect 78728 35416 79001 35428
rect 80510 35416 81015 36141
rect 100968 36307 101045 36361
rect 100968 36103 101046 36307
rect 103010 36203 103515 36368
rect 123260 36342 123795 37061
rect 101149 36183 103515 36203
rect 101149 36150 101157 36183
rect 101191 36150 103515 36183
rect 101149 36141 103515 36150
rect 100968 35428 100974 36103
rect 101038 35428 101046 36103
rect 100968 35419 101046 35428
rect 101076 36103 101154 36113
rect 101076 35428 101083 36103
rect 101147 35428 101154 36103
rect 101076 35416 101154 35428
rect 101278 36103 101366 36114
rect 101278 35428 101284 36103
rect 101359 35842 101366 36103
rect 101359 35428 101569 35842
rect 101278 35416 101569 35428
rect 103010 35416 103515 36141
rect 123468 36307 123545 36342
rect 123468 36103 123546 36307
rect 125510 36203 126015 36368
rect 145815 36356 146238 36779
rect 123649 36183 126015 36203
rect 123649 36150 123657 36183
rect 123649 36149 123691 36150
rect 123860 36149 126015 36183
rect 123649 36141 126015 36149
rect 125242 36140 126015 36141
rect 123468 35428 123474 36103
rect 123538 35428 123546 36103
rect 123576 36103 123654 36113
rect 123576 35605 123583 36103
rect 123468 35419 123546 35428
rect 123573 35428 123583 35605
rect 123647 35428 123654 36103
rect 123573 35416 123654 35428
rect 123878 36103 123966 36114
rect 123878 35428 123884 36103
rect 123959 36098 123966 36103
rect 123959 35741 123971 36098
rect 123959 35428 124041 35741
rect 123878 35416 124041 35428
rect 125510 35416 126015 36140
rect 145968 36307 146045 36356
rect 145968 36103 146046 36307
rect 148010 36203 148515 36368
rect 146149 36183 148515 36203
rect 146149 36150 146157 36183
rect 146149 36148 146178 36150
rect 146552 36148 148515 36183
rect 146149 36141 148515 36148
rect 145968 35428 145974 36103
rect 146038 35428 146046 36103
rect 145968 35419 146046 35428
rect 146076 36103 146154 36113
rect 146076 35428 146083 36103
rect 146147 35428 146154 36103
rect 146076 35416 146154 35428
rect 146574 36103 146708 36114
rect 146574 35428 146584 36103
rect 146659 35946 146708 36103
rect 146659 35428 146737 35946
rect 56074 35201 56131 35416
rect 53981 35083 56131 35201
rect 53981 34470 56124 35083
rect 56225 34732 56618 35416
rect 78575 35039 78651 35416
rect 76485 34732 78651 35039
rect 78757 34732 79001 35416
rect 101081 35072 101147 35416
rect 98992 34998 101147 35072
rect 98992 34732 101136 34998
rect 101291 34732 101569 35416
rect 123573 35008 123651 35416
rect 121580 34732 123651 35008
rect 123890 34732 124041 35416
rect 146077 35011 146141 35416
rect 146574 35399 146737 35428
rect 148010 35416 148515 36141
rect 146593 35280 146737 35399
rect 53983 34250 54481 34470
rect 56225 34426 56691 34732
rect 53980 32650 54485 34250
rect 56256 33053 56691 34426
rect 76480 34645 78651 34732
rect 76480 34339 78634 34645
rect 76480 34242 76989 34339
rect 56172 32078 56822 33053
rect 76480 32650 76985 34242
rect 78756 33205 79191 34732
rect 98977 34613 101136 34732
rect 98977 34250 99481 34613
rect 98977 34223 99485 34250
rect 78639 32054 79419 33205
rect 98980 32650 99485 34223
rect 101256 33010 101691 34732
rect 101237 32650 101691 33010
rect 121480 34709 123651 34732
rect 121480 34237 123632 34709
rect 121480 32650 121985 34237
rect 123864 34171 124191 34732
rect 143962 34194 146141 35011
rect 146575 34740 147175 35280
rect 146550 34350 147175 34740
rect 123756 32981 124191 34171
rect 123746 32846 124281 32981
rect 123738 32650 124281 32846
rect 143980 32650 144485 34194
rect 146550 34005 147150 34350
rect 146415 33810 147150 34005
rect 146415 33644 147015 33810
rect 146256 33490 147015 33644
rect 146256 33060 147265 33490
rect 146238 33015 147265 33060
rect 101237 32113 101683 32650
rect 123746 32262 124281 32650
rect 146238 32125 147295 33015
rect 146695 32085 147295 32125
rect 55624 13329 56240 13843
rect 55958 13103 56036 13329
rect 58010 13204 58515 13368
rect 77978 13353 78742 13800
rect 57750 13203 58515 13204
rect 56139 13183 58515 13203
rect 56139 13150 56147 13183
rect 56191 13150 58515 13183
rect 56139 13141 58515 13150
rect 53915 3032 54493 10407
rect 55958 3128 55964 13103
rect 56028 3128 56036 13103
rect 55958 3119 56036 3128
rect 56066 13103 56144 13113
rect 56066 3128 56073 13103
rect 56137 3128 56144 13103
rect 56066 3032 56144 3128
rect 56203 13103 56291 13114
rect 56203 3128 56209 13103
rect 56284 3128 56291 13103
rect 58010 12539 58515 13141
rect 78468 13307 78545 13353
rect 78468 13103 78546 13307
rect 80510 13203 81015 13368
rect 100593 13341 101248 13949
rect 78649 13183 81015 13203
rect 78649 13150 78657 13183
rect 78691 13150 81015 13183
rect 78649 13141 81015 13150
rect 56203 3116 56291 3128
rect 76608 3078 76986 10846
rect 78468 3128 78474 13103
rect 78538 3128 78546 13103
rect 78468 3119 78546 3128
rect 78576 13103 78654 13113
rect 78576 3128 78583 13103
rect 78647 3128 78654 13103
rect 78576 3078 78654 3128
rect 78728 13103 78816 13114
rect 78728 3128 78734 13103
rect 78809 3128 78816 13103
rect 80510 12585 81015 13141
rect 100968 13307 101045 13341
rect 100968 13103 101046 13307
rect 103010 13203 103515 13368
rect 122926 13359 123745 13810
rect 101149 13183 103515 13203
rect 101149 13150 101157 13183
rect 101191 13150 103515 13183
rect 101149 13141 103515 13150
rect 78728 3116 78816 3128
rect 53915 2661 56146 3032
rect 76608 3009 78654 3078
rect 98931 3028 99491 10748
rect 100968 3128 100974 13103
rect 101038 3128 101046 13103
rect 100968 3119 101046 3128
rect 101076 13103 101154 13113
rect 101076 3128 101083 13103
rect 101147 3128 101154 13103
rect 101076 3028 101154 3128
rect 101278 13103 101366 13114
rect 101278 3128 101284 13103
rect 101359 3128 101366 13103
rect 103010 12713 103515 13141
rect 123468 13307 123545 13359
rect 123468 13103 123546 13307
rect 125510 13203 126015 13368
rect 145461 13361 146244 13652
rect 123649 13183 126015 13203
rect 123649 13150 123657 13183
rect 123649 13149 123691 13150
rect 123860 13149 126015 13183
rect 123649 13141 126015 13149
rect 125242 13140 126015 13141
rect 101278 3116 101366 3128
rect 76608 2644 78651 3009
rect 98931 2608 101154 3028
rect 121419 3037 121964 10751
rect 123468 3128 123474 13103
rect 123538 3128 123546 13103
rect 123468 3119 123546 3128
rect 123576 13103 123654 13113
rect 123576 3128 123583 13103
rect 123647 3128 123654 13103
rect 123576 3037 123654 3128
rect 123878 13103 123966 13114
rect 123878 3128 123884 13103
rect 123959 13098 123966 13103
rect 123959 13077 123971 13098
rect 123959 3128 124014 13077
rect 125510 12199 126015 13140
rect 145968 13307 146045 13361
rect 145968 13103 146046 13307
rect 148010 13203 148515 13368
rect 146149 13183 148515 13203
rect 146149 13150 146157 13183
rect 146149 13148 146178 13150
rect 146552 13148 148515 13183
rect 146149 13141 148515 13148
rect 146578 13113 146666 13114
rect 123878 3116 124014 3128
rect 123931 3082 124014 3116
rect 121419 2979 123654 3037
rect 143922 3072 144486 10752
rect 145968 3128 145974 13103
rect 146038 3128 146046 13103
rect 145968 3119 146046 3128
rect 146076 13103 146154 13113
rect 146076 3128 146083 13103
rect 146147 3128 146154 13103
rect 146076 3072 146154 3128
rect 121419 2592 123650 2979
rect 143922 2974 146154 3072
rect 146564 13103 146691 13113
rect 146564 3128 146584 13103
rect 146659 3128 146691 13103
rect 148010 12577 148515 13141
rect 146564 3040 146691 3128
rect 143922 2641 146149 2974
use BarePadArray1x5  BarePadArray1x5_0
timestamp 1663655995
transform 1 0 44875 0 1 695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_1
timestamp 1663655995
transform 1 0 44875 0 1 23695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_2
timestamp 1663655995
transform 1 0 44875 0 1 46695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_3
timestamp 1663655995
transform 1 0 44875 0 1 69695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_4
timestamp 1663655995
transform 1 0 44875 0 1 92695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_5
timestamp 1663655995
transform 1 0 44875 0 1 115695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_6
timestamp 1663655995
transform 1 0 44875 0 1 138695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_7
timestamp 1663655995
transform 1 0 44875 0 1 161695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_8
timestamp 1663655995
transform 1 0 44875 0 1 184695
box 115 -840 112615 22160
use BarePadArray1x5  BarePadArray1x5_9
timestamp 1663655995
transform 1 0 44875 0 1 207695
box 115 -840 112615 22160
<< end >>
