magic
tech sky130A
timestamp 1663612738
<< nwell >>
rect 1295 -920 3620 -620
rect 2445 -1130 3620 -920
<< pwell >>
rect 1130 -1125 2395 -1010
rect 1125 -1170 2395 -1125
rect 1130 -1230 2395 -1170
rect 1125 -1275 2395 -1230
rect 1130 -1330 2395 -1275
rect 2520 -1305 2675 -1265
rect 2945 -1305 3005 -1265
rect 1130 -1360 3620 -1330
rect 1125 -1400 3620 -1360
rect 1130 -1410 3620 -1400
rect 1125 -1455 3620 -1410
rect 1130 -1835 3620 -1455
<< pmoslvt >>
rect 1415 -870 1515 -670
rect 1615 -870 1715 -670
rect 2540 -1070 2590 -670
rect 2820 -1070 2870 -670
rect 3105 -1070 3155 -670
rect 3390 -1070 3440 -670
<< nmoslvt >>
rect 1560 -1295 1610 -1195
rect 1660 -1295 1710 -1195
rect 2160 -1240 2210 -1040
rect 2260 -1240 2310 -1040
rect 1285 -1770 1385 -1470
rect 1485 -1770 1585 -1470
rect 1885 -1770 1985 -1470
rect 2085 -1770 2185 -1470
rect 2485 -1770 2585 -1470
rect 2820 -1670 2870 -1470
rect 3105 -1670 3155 -1470
rect 3390 -1670 3440 -1470
<< ndiff >>
rect 2110 -1050 2160 -1040
rect 1510 -1205 1560 -1195
rect 1510 -1280 1525 -1205
rect 1545 -1280 1560 -1205
rect 1510 -1295 1560 -1280
rect 1610 -1205 1660 -1195
rect 1610 -1280 1625 -1205
rect 1645 -1280 1660 -1205
rect 1610 -1295 1660 -1280
rect 1710 -1205 1760 -1195
rect 1710 -1280 1725 -1205
rect 1745 -1280 1760 -1205
rect 2110 -1230 2120 -1050
rect 2150 -1230 2160 -1050
rect 2110 -1240 2160 -1230
rect 2210 -1050 2260 -1040
rect 2210 -1230 2220 -1050
rect 2250 -1230 2260 -1050
rect 2210 -1240 2260 -1230
rect 2310 -1050 2360 -1040
rect 2310 -1230 2320 -1050
rect 2350 -1230 2360 -1050
rect 2310 -1240 2360 -1230
rect 1710 -1295 1760 -1280
rect 1185 -1495 1285 -1470
rect 1185 -1750 1205 -1495
rect 1265 -1750 1285 -1495
rect 1185 -1770 1285 -1750
rect 1385 -1495 1485 -1470
rect 1385 -1750 1405 -1495
rect 1465 -1750 1485 -1495
rect 1385 -1770 1485 -1750
rect 1585 -1495 1685 -1470
rect 1785 -1495 1885 -1470
rect 1585 -1750 1605 -1495
rect 1665 -1750 1685 -1495
rect 1785 -1750 1805 -1495
rect 1865 -1750 1885 -1495
rect 1585 -1770 1685 -1750
rect 1785 -1770 1885 -1750
rect 1985 -1495 2085 -1470
rect 1985 -1750 2005 -1495
rect 2065 -1750 2085 -1495
rect 1985 -1770 2085 -1750
rect 2185 -1495 2285 -1470
rect 2385 -1495 2485 -1470
rect 2185 -1750 2205 -1495
rect 2265 -1750 2285 -1495
rect 2385 -1750 2405 -1495
rect 2465 -1750 2485 -1495
rect 2185 -1770 2285 -1750
rect 2385 -1770 2485 -1750
rect 2585 -1495 2685 -1470
rect 2585 -1750 2605 -1495
rect 2665 -1750 2685 -1495
rect 2750 -1485 2820 -1470
rect 2750 -1655 2765 -1485
rect 2805 -1655 2820 -1485
rect 2750 -1670 2820 -1655
rect 2870 -1485 2940 -1470
rect 2870 -1655 2885 -1485
rect 2925 -1655 2940 -1485
rect 2870 -1670 2940 -1655
rect 3035 -1485 3105 -1470
rect 3035 -1655 3050 -1485
rect 3090 -1655 3105 -1485
rect 3035 -1670 3105 -1655
rect 3155 -1485 3225 -1470
rect 3155 -1655 3170 -1485
rect 3210 -1655 3225 -1485
rect 3155 -1670 3225 -1655
rect 3320 -1485 3390 -1470
rect 3320 -1655 3335 -1485
rect 3375 -1655 3390 -1485
rect 3320 -1670 3390 -1655
rect 3440 -1485 3510 -1470
rect 3440 -1655 3455 -1485
rect 3495 -1655 3510 -1485
rect 3440 -1670 3510 -1655
rect 2585 -1770 2685 -1750
<< pdiff >>
rect 1315 -690 1415 -670
rect 1315 -850 1335 -690
rect 1395 -850 1415 -690
rect 1315 -870 1415 -850
rect 1515 -690 1615 -670
rect 1515 -850 1535 -690
rect 1595 -850 1615 -690
rect 1515 -870 1615 -850
rect 1715 -690 1815 -670
rect 1715 -850 1735 -690
rect 1795 -850 1815 -690
rect 1715 -870 1815 -850
rect 2470 -685 2540 -670
rect 2470 -1055 2485 -685
rect 2525 -1055 2540 -685
rect 2470 -1070 2540 -1055
rect 2590 -685 2660 -670
rect 2745 -685 2820 -670
rect 2590 -1055 2605 -685
rect 2645 -1055 2660 -685
rect 2745 -1055 2765 -685
rect 2805 -1055 2820 -685
rect 2590 -1070 2660 -1055
rect 2745 -1070 2820 -1055
rect 2870 -685 2940 -670
rect 3030 -685 3105 -670
rect 2870 -1055 2885 -685
rect 2925 -1055 2940 -685
rect 3030 -1055 3050 -685
rect 3090 -1055 3105 -685
rect 2870 -1070 2940 -1055
rect 3030 -1070 3105 -1055
rect 3155 -685 3225 -670
rect 3315 -685 3390 -670
rect 3155 -1055 3170 -685
rect 3210 -1055 3225 -685
rect 3315 -1055 3335 -685
rect 3375 -1055 3390 -685
rect 3155 -1070 3225 -1055
rect 3315 -1070 3390 -1055
rect 3440 -685 3510 -670
rect 3440 -1055 3455 -685
rect 3495 -1055 3510 -685
rect 3440 -1070 3510 -1055
<< ndiffc >>
rect 1525 -1280 1545 -1205
rect 1625 -1280 1645 -1205
rect 1725 -1280 1745 -1205
rect 2120 -1230 2150 -1050
rect 2220 -1230 2250 -1050
rect 2320 -1230 2350 -1050
rect 1205 -1750 1265 -1495
rect 1405 -1750 1465 -1495
rect 1605 -1750 1665 -1495
rect 1805 -1750 1865 -1495
rect 2005 -1750 2065 -1495
rect 2205 -1750 2265 -1495
rect 2405 -1750 2465 -1495
rect 2605 -1750 2665 -1495
rect 2765 -1655 2805 -1485
rect 2885 -1655 2925 -1485
rect 3050 -1655 3090 -1485
rect 3170 -1655 3210 -1485
rect 3335 -1655 3375 -1485
rect 3455 -1655 3495 -1485
<< pdiffc >>
rect 1335 -850 1395 -690
rect 1535 -850 1595 -690
rect 1735 -850 1795 -690
rect 2485 -1055 2525 -685
rect 2605 -1055 2645 -685
rect 2765 -1055 2805 -685
rect 2885 -1055 2925 -685
rect 3050 -1055 3090 -685
rect 3170 -1055 3210 -685
rect 3335 -1055 3375 -685
rect 3455 -1055 3495 -685
<< psubdiff >>
rect 1685 -1495 1785 -1470
rect 1685 -1750 1705 -1495
rect 1765 -1750 1785 -1495
rect 1685 -1770 1785 -1750
rect 2285 -1495 2385 -1470
rect 2285 -1750 2305 -1495
rect 2365 -1750 2385 -1495
rect 2285 -1770 2385 -1750
rect 2940 -1480 3035 -1470
rect 2940 -1660 2965 -1480
rect 3005 -1660 3035 -1480
rect 2940 -1670 3035 -1660
rect 3225 -1480 3320 -1470
rect 3225 -1660 3250 -1480
rect 3290 -1660 3320 -1480
rect 3225 -1670 3320 -1660
rect 3510 -1480 3595 -1470
rect 3510 -1660 3535 -1480
rect 3575 -1660 3595 -1480
rect 3510 -1670 3595 -1660
<< nsubdiff >>
rect 1815 -690 1915 -670
rect 1815 -850 1840 -690
rect 1895 -850 1915 -690
rect 1815 -870 1915 -850
rect 2660 -685 2745 -670
rect 2660 -1055 2685 -685
rect 2725 -1055 2745 -685
rect 2660 -1070 2745 -1055
rect 2940 -685 3030 -670
rect 2940 -1055 2965 -685
rect 3005 -1055 3030 -685
rect 2940 -1070 3030 -1055
rect 3225 -685 3315 -670
rect 3225 -1055 3250 -685
rect 3290 -1055 3315 -685
rect 3225 -1070 3315 -1055
rect 3510 -685 3595 -670
rect 3510 -1055 3535 -685
rect 3575 -1055 3595 -685
rect 3510 -1070 3595 -1055
<< psubdiffcont >>
rect 1705 -1750 1765 -1495
rect 2305 -1750 2365 -1495
rect 2965 -1660 3005 -1480
rect 3250 -1660 3290 -1480
rect 3535 -1660 3575 -1480
<< nsubdiffcont >>
rect 1840 -850 1895 -690
rect 2685 -1055 2725 -685
rect 2965 -1055 3005 -685
rect 3250 -1055 3290 -685
rect 3535 -1055 3575 -685
<< poly >>
rect 1415 -670 1515 -635
rect 1615 -670 1715 -635
rect 2540 -670 2590 -650
rect 2820 -670 2870 -650
rect 3105 -670 3155 -650
rect 3390 -670 3440 -650
rect 1415 -895 1515 -870
rect 1415 -935 1425 -895
rect 1505 -900 1515 -895
rect 1615 -900 1715 -870
rect 1505 -935 1715 -900
rect 1415 -945 1715 -935
rect 2160 -1040 2210 -1015
rect 2260 -1040 2310 -1015
rect 1645 -1145 1710 -1135
rect 1645 -1165 1655 -1145
rect 1700 -1165 1710 -1145
rect 1645 -1175 1710 -1165
rect 1560 -1195 1610 -1175
rect 1660 -1195 1710 -1175
rect 2540 -1095 2590 -1070
rect 2540 -1115 2545 -1095
rect 2580 -1115 2590 -1095
rect 2540 -1125 2590 -1115
rect 2820 -1135 2870 -1070
rect 3105 -1135 3155 -1070
rect 3390 -1135 3440 -1070
rect 2780 -1145 2870 -1135
rect 2780 -1175 2790 -1145
rect 2860 -1175 2870 -1145
rect 2780 -1185 2870 -1175
rect 3065 -1145 3155 -1135
rect 3065 -1175 3075 -1145
rect 3145 -1175 3155 -1145
rect 3065 -1185 3155 -1175
rect 3350 -1145 3440 -1135
rect 3350 -1175 3360 -1145
rect 3430 -1175 3440 -1145
rect 3350 -1185 3440 -1175
rect 2160 -1265 2210 -1240
rect 2145 -1275 2210 -1265
rect 1560 -1310 1610 -1295
rect 1660 -1310 1710 -1295
rect 2145 -1310 2155 -1275
rect 2185 -1310 2210 -1275
rect 1530 -1320 1610 -1310
rect 2145 -1320 2210 -1310
rect 2260 -1265 2310 -1240
rect 2260 -1275 2325 -1265
rect 2260 -1310 2285 -1275
rect 2315 -1310 2325 -1275
rect 2260 -1320 2325 -1310
rect 1530 -1340 1540 -1320
rect 1585 -1340 1610 -1320
rect 1530 -1350 1610 -1340
rect 1885 -1355 1980 -1340
rect 1885 -1390 1895 -1355
rect 1970 -1390 1980 -1355
rect 1885 -1410 1980 -1390
rect 2485 -1405 2585 -1395
rect 1285 -1415 1585 -1410
rect 1285 -1450 1295 -1415
rect 1370 -1450 1585 -1415
rect 1285 -1460 1585 -1450
rect 1285 -1470 1385 -1460
rect 1485 -1470 1585 -1460
rect 1885 -1460 2185 -1410
rect 1885 -1470 1985 -1460
rect 2085 -1470 2185 -1460
rect 2485 -1440 2500 -1405
rect 2575 -1440 2585 -1405
rect 2485 -1470 2585 -1440
rect 2820 -1470 2870 -1185
rect 3105 -1470 3155 -1185
rect 3390 -1470 3440 -1185
rect 2820 -1685 2870 -1670
rect 3105 -1685 3155 -1670
rect 3390 -1685 3440 -1670
rect 1285 -1805 1385 -1770
rect 1485 -1805 1585 -1770
rect 1885 -1805 1985 -1770
rect 2085 -1805 2185 -1770
rect 2485 -1805 2585 -1770
<< polycont >>
rect 1425 -935 1505 -895
rect 1655 -1165 1700 -1145
rect 2545 -1115 2580 -1095
rect 2790 -1175 2860 -1145
rect 3075 -1175 3145 -1145
rect 3360 -1175 3430 -1145
rect 2155 -1310 2185 -1275
rect 2285 -1310 2315 -1275
rect 1540 -1340 1585 -1320
rect 1895 -1390 1970 -1355
rect 1295 -1450 1370 -1415
rect 2500 -1440 2575 -1405
<< locali >>
rect 1325 -690 1405 -680
rect 1325 -850 1335 -690
rect 1395 -850 1405 -690
rect 1325 -860 1405 -850
rect 1525 -690 1605 -680
rect 1525 -850 1535 -690
rect 1595 -850 1605 -690
rect 1525 -860 1605 -850
rect 1725 -690 1805 -680
rect 1725 -850 1735 -690
rect 1795 -850 1805 -690
rect 1725 -860 1805 -850
rect 1830 -690 1905 -680
rect 1830 -850 1840 -690
rect 1895 -850 1905 -690
rect 1830 -860 1905 -850
rect 2475 -685 2535 -675
rect 1325 -895 1395 -860
rect 1415 -895 1515 -875
rect 1325 -935 1425 -895
rect 1505 -935 1515 -895
rect 1325 -945 1515 -935
rect 2315 -920 2440 -915
rect 1325 -950 1415 -945
rect 2315 -955 2325 -920
rect 2345 -955 2440 -920
rect 2315 -965 2440 -955
rect 2115 -1050 2155 -1040
rect 2115 -1080 2120 -1050
rect 1510 -1085 2120 -1080
rect 1510 -1105 1515 -1085
rect 1545 -1105 2120 -1085
rect 1510 -1110 2120 -1105
rect 1445 -1140 1710 -1135
rect 1445 -1160 1450 -1140
rect 1480 -1145 1710 -1140
rect 1480 -1160 1655 -1145
rect 1445 -1165 1655 -1160
rect 1700 -1165 1710 -1145
rect 1645 -1175 1710 -1165
rect 1510 -1205 1555 -1195
rect 1510 -1280 1520 -1205
rect 1545 -1280 1555 -1205
rect 1510 -1290 1555 -1280
rect 1615 -1205 1655 -1195
rect 1615 -1280 1625 -1205
rect 1645 -1280 1655 -1205
rect 1530 -1320 1595 -1310
rect 1530 -1340 1540 -1320
rect 1585 -1340 1595 -1320
rect 1530 -1350 1595 -1340
rect 1195 -1415 1475 -1410
rect 1195 -1450 1295 -1415
rect 1370 -1450 1475 -1415
rect 1195 -1460 1475 -1450
rect 1195 -1495 1275 -1460
rect 1615 -1485 1655 -1280
rect 1715 -1205 1760 -1195
rect 1715 -1280 1725 -1205
rect 1750 -1280 1760 -1205
rect 2115 -1230 2120 -1110
rect 2150 -1230 2155 -1050
rect 2115 -1240 2155 -1230
rect 2215 -1050 2255 -1040
rect 2215 -1230 2220 -1050
rect 2250 -1230 2255 -1050
rect 1715 -1290 1760 -1280
rect 2145 -1275 2195 -1265
rect 1890 -1355 1975 -1345
rect 1890 -1390 1895 -1355
rect 1970 -1390 1975 -1355
rect 2145 -1350 2155 -1275
rect 2185 -1350 2195 -1275
rect 2145 -1385 2195 -1350
rect 1890 -1415 1975 -1390
rect 1795 -1455 2075 -1415
rect 1195 -1750 1205 -1495
rect 1265 -1750 1275 -1495
rect 1195 -1760 1275 -1750
rect 1395 -1495 1475 -1485
rect 1395 -1750 1405 -1495
rect 1465 -1750 1475 -1495
rect 1395 -1760 1475 -1750
rect 1595 -1495 1675 -1485
rect 1595 -1750 1605 -1495
rect 1665 -1750 1675 -1495
rect 1595 -1760 1675 -1750
rect 1695 -1495 1775 -1480
rect 1695 -1750 1705 -1495
rect 1765 -1750 1775 -1495
rect 1695 -1760 1775 -1750
rect 1795 -1495 1875 -1455
rect 2215 -1485 2255 -1230
rect 2315 -1050 2355 -965
rect 2315 -1230 2320 -1050
rect 2350 -1230 2355 -1050
rect 2400 -1085 2440 -965
rect 2475 -1055 2485 -685
rect 2525 -1055 2535 -685
rect 2475 -1065 2535 -1055
rect 2595 -685 2655 -675
rect 2595 -1055 2605 -685
rect 2645 -1055 2655 -685
rect 2595 -1065 2655 -1055
rect 2675 -685 2735 -675
rect 2675 -1055 2685 -685
rect 2725 -1055 2735 -685
rect 2675 -1065 2735 -1055
rect 2755 -685 2815 -675
rect 2755 -1055 2765 -685
rect 2805 -1055 2815 -685
rect 2755 -1065 2815 -1055
rect 2875 -685 2935 -675
rect 2875 -1055 2885 -685
rect 2925 -1055 2935 -685
rect 2875 -1065 2935 -1055
rect 2955 -685 3015 -675
rect 2955 -1055 2965 -685
rect 3005 -1055 3015 -685
rect 2955 -1065 3015 -1055
rect 3040 -685 3100 -675
rect 3040 -1055 3050 -685
rect 3090 -1055 3100 -685
rect 3040 -1065 3100 -1055
rect 3160 -685 3220 -675
rect 3160 -1055 3170 -685
rect 3210 -1055 3220 -685
rect 3160 -1065 3220 -1055
rect 3240 -685 3300 -675
rect 3240 -1055 3250 -685
rect 3290 -1055 3300 -685
rect 3240 -1065 3300 -1055
rect 3325 -685 3385 -675
rect 3325 -1055 3335 -685
rect 3375 -1055 3385 -685
rect 3325 -1065 3385 -1055
rect 3445 -685 3505 -675
rect 3445 -1055 3455 -685
rect 3495 -1055 3505 -685
rect 3445 -1065 3505 -1055
rect 3525 -685 3585 -675
rect 3525 -1055 3535 -685
rect 3575 -1055 3585 -685
rect 3525 -1065 3585 -1055
rect 2400 -1095 2590 -1085
rect 2400 -1115 2545 -1095
rect 2580 -1115 2590 -1095
rect 2400 -1125 2590 -1115
rect 2780 -1145 2870 -1135
rect 2780 -1175 2790 -1145
rect 2860 -1175 2870 -1145
rect 2780 -1185 2870 -1175
rect 3065 -1145 3155 -1135
rect 3065 -1175 3075 -1145
rect 3145 -1175 3155 -1145
rect 3065 -1185 3155 -1175
rect 3350 -1145 3440 -1135
rect 3350 -1175 3360 -1145
rect 3430 -1175 3440 -1145
rect 3350 -1185 3440 -1175
rect 2315 -1240 2355 -1230
rect 2275 -1275 2325 -1265
rect 2520 -1275 3005 -1265
rect 2275 -1310 2285 -1275
rect 2520 -1295 2530 -1275
rect 2570 -1295 2955 -1275
rect 2995 -1295 3005 -1275
rect 2315 -1310 2325 -1300
rect 2520 -1305 3005 -1295
rect 2275 -1320 2325 -1310
rect 2520 -1345 2735 -1335
rect 2520 -1365 2530 -1345
rect 2570 -1365 2685 -1345
rect 2725 -1365 2735 -1345
rect 2520 -1375 2735 -1365
rect 2485 -1405 2585 -1395
rect 2485 -1440 2500 -1405
rect 2575 -1440 2585 -1405
rect 2485 -1455 2585 -1440
rect 1795 -1750 1805 -1495
rect 1865 -1750 1875 -1495
rect 1795 -1760 1875 -1750
rect 1995 -1495 2075 -1485
rect 1995 -1750 2005 -1495
rect 2065 -1750 2075 -1495
rect 1995 -1760 2075 -1750
rect 2195 -1495 2275 -1485
rect 2195 -1750 2205 -1495
rect 2265 -1750 2275 -1495
rect 2195 -1760 2275 -1750
rect 2295 -1495 2375 -1480
rect 2295 -1750 2305 -1495
rect 2365 -1750 2375 -1495
rect 2295 -1760 2375 -1750
rect 2395 -1495 2475 -1480
rect 2395 -1750 2405 -1495
rect 2465 -1750 2475 -1495
rect 2395 -1760 2475 -1750
rect 2595 -1495 2675 -1480
rect 2595 -1750 2605 -1495
rect 2665 -1750 2675 -1495
rect 2755 -1485 2815 -1475
rect 2755 -1655 2765 -1485
rect 2805 -1655 2815 -1485
rect 2755 -1665 2815 -1655
rect 2875 -1485 2935 -1475
rect 2875 -1655 2885 -1485
rect 2925 -1655 2935 -1485
rect 2875 -1665 2935 -1655
rect 2955 -1480 3015 -1475
rect 2955 -1660 2965 -1480
rect 3005 -1660 3015 -1480
rect 2955 -1665 3015 -1660
rect 3040 -1485 3100 -1475
rect 3040 -1655 3050 -1485
rect 3090 -1655 3100 -1485
rect 3040 -1665 3100 -1655
rect 3160 -1485 3220 -1475
rect 3160 -1655 3170 -1485
rect 3210 -1655 3220 -1485
rect 3160 -1665 3220 -1655
rect 3240 -1480 3300 -1475
rect 3240 -1660 3250 -1480
rect 3290 -1660 3300 -1480
rect 3240 -1665 3300 -1660
rect 3325 -1485 3385 -1475
rect 3325 -1655 3335 -1485
rect 3375 -1655 3385 -1485
rect 3325 -1665 3385 -1655
rect 3445 -1485 3505 -1475
rect 3445 -1655 3455 -1485
rect 3495 -1655 3505 -1485
rect 3445 -1665 3505 -1655
rect 3525 -1480 3585 -1475
rect 3525 -1660 3535 -1480
rect 3575 -1660 3585 -1480
rect 3525 -1665 3585 -1660
rect 2595 -1760 2675 -1750
<< viali >>
rect 1340 -845 1390 -695
rect 1540 -845 1590 -695
rect 1740 -845 1790 -695
rect 1840 -850 1895 -690
rect 1425 -935 1505 -895
rect 2325 -955 2345 -920
rect 1515 -1105 1545 -1085
rect 1450 -1160 1480 -1140
rect 1520 -1280 1525 -1205
rect 1525 -1280 1540 -1205
rect 1540 -1340 1585 -1320
rect 1300 -1445 1365 -1420
rect 1730 -1280 1745 -1205
rect 1745 -1280 1750 -1205
rect 1900 -1385 1965 -1360
rect 2155 -1310 2185 -1295
rect 2155 -1350 2185 -1310
rect 1405 -1750 1465 -1495
rect 1705 -1750 1765 -1495
rect 2485 -1055 2525 -685
rect 2610 -1045 2640 -695
rect 2685 -1055 2725 -685
rect 2765 -1055 2805 -685
rect 2890 -1045 2920 -695
rect 2965 -1055 3005 -685
rect 3050 -1055 3090 -685
rect 3175 -1045 3205 -695
rect 3250 -1055 3290 -685
rect 3335 -1055 3375 -685
rect 3460 -1045 3490 -695
rect 3535 -1055 3575 -685
rect 2790 -1175 2860 -1145
rect 3075 -1175 3145 -1145
rect 3360 -1175 3430 -1145
rect 2285 -1300 2315 -1275
rect 2315 -1300 2335 -1275
rect 2530 -1295 2570 -1275
rect 2955 -1295 2995 -1275
rect 2530 -1365 2570 -1345
rect 2685 -1365 2725 -1345
rect 2505 -1435 2570 -1410
rect 2005 -1750 2065 -1495
rect 2305 -1750 2365 -1495
rect 2405 -1750 2465 -1495
rect 2610 -1745 2660 -1500
rect 2770 -1645 2800 -1495
rect 2890 -1645 2920 -1495
rect 2970 -1645 3000 -1495
rect 3055 -1648 3085 -1498
rect 3175 -1645 3205 -1495
rect 3255 -1641 3285 -1491
rect 3339 -1646 3369 -1496
rect 3460 -1645 3490 -1495
rect 3541 -1643 3571 -1493
<< metal1 >>
rect 1200 40 3585 90
rect 1200 -5 1255 40
rect 1305 -5 1355 40
rect 1405 -5 1455 40
rect 1505 -5 1555 40
rect 1605 -5 1655 40
rect 1705 -5 1755 40
rect 1805 -5 1855 40
rect 1905 -5 1955 40
rect 2005 -5 2055 40
rect 2105 -5 2155 40
rect 2205 -5 2255 40
rect 2305 -5 2355 40
rect 2405 -5 2455 40
rect 2505 -5 2555 40
rect 2605 -5 2655 40
rect 2705 -5 2755 40
rect 2805 -5 2855 40
rect 2905 -5 2955 40
rect 3005 -5 3055 40
rect 3105 -5 3155 40
rect 3205 -5 3255 40
rect 3305 -5 3355 40
rect 3405 -5 3455 40
rect 3505 -5 3585 40
rect 1200 -35 3585 -5
rect 1200 -80 1255 -35
rect 1305 -80 1355 -35
rect 1405 -80 1455 -35
rect 1505 -80 1555 -35
rect 1605 -80 1655 -35
rect 1705 -80 1755 -35
rect 1805 -80 1855 -35
rect 1905 -80 1955 -35
rect 2005 -80 2055 -35
rect 2105 -80 2155 -35
rect 2205 -80 2255 -35
rect 2305 -80 2355 -35
rect 2405 -80 2455 -35
rect 2505 -80 2555 -35
rect 2605 -80 2655 -35
rect 2705 -80 2755 -35
rect 2805 -80 2855 -35
rect 2905 -80 2955 -35
rect 3005 -80 3055 -35
rect 3105 -80 3155 -35
rect 3205 -80 3255 -35
rect 3305 -80 3355 -35
rect 3405 -80 3455 -35
rect 3505 -80 3585 -35
rect 1200 -110 3585 -80
rect 1200 -155 1255 -110
rect 1305 -155 1355 -110
rect 1405 -155 1455 -110
rect 1505 -155 1555 -110
rect 1605 -155 1655 -110
rect 1705 -155 1755 -110
rect 1805 -155 1855 -110
rect 1905 -155 1955 -110
rect 2005 -155 2055 -110
rect 2105 -155 2155 -110
rect 2205 -155 2255 -110
rect 2305 -155 2355 -110
rect 2405 -155 2455 -110
rect 2505 -155 2555 -110
rect 2605 -155 2655 -110
rect 2705 -155 2755 -110
rect 2805 -155 2855 -110
rect 2905 -155 2955 -110
rect 3005 -155 3055 -110
rect 3105 -155 3155 -110
rect 3205 -155 3255 -110
rect 3305 -155 3355 -110
rect 3405 -155 3455 -110
rect 3505 -155 3585 -110
rect 1200 -560 3585 -155
rect 1125 -620 3620 -560
rect 1330 -695 1400 -685
rect 1330 -845 1340 -695
rect 1390 -845 1400 -695
rect 1330 -895 1400 -845
rect 1530 -695 1600 -620
rect 1530 -845 1540 -695
rect 1590 -845 1600 -695
rect 1530 -855 1600 -845
rect 1730 -695 1800 -685
rect 1730 -845 1740 -695
rect 1790 -845 1800 -695
rect 1415 -895 1515 -880
rect 1325 -935 1425 -895
rect 1505 -935 1515 -895
rect 1325 -945 1515 -935
rect 1430 -1000 1515 -945
rect 1730 -915 1800 -845
rect 1830 -690 1905 -620
rect 1830 -850 1840 -690
rect 1895 -850 1905 -690
rect 1830 -860 1905 -850
rect 2475 -685 2535 -620
rect 1730 -920 2355 -915
rect 1730 -955 2325 -920
rect 2345 -955 2355 -920
rect 1730 -965 2355 -955
rect 1430 -1035 1550 -1000
rect 1730 -1015 1800 -965
rect 1510 -1085 1550 -1035
rect 1510 -1105 1515 -1085
rect 1545 -1105 1550 -1085
rect 1125 -1140 1485 -1125
rect 1125 -1160 1450 -1140
rect 1480 -1160 1485 -1140
rect 1125 -1170 1485 -1160
rect 1510 -1205 1550 -1105
rect 1125 -1275 1480 -1230
rect 1435 -1310 1480 -1275
rect 1510 -1280 1520 -1205
rect 1540 -1280 1550 -1205
rect 1510 -1285 1550 -1280
rect 1720 -1050 1800 -1015
rect 1720 -1205 1760 -1050
rect 2475 -1055 2485 -685
rect 2525 -1055 2535 -685
rect 2475 -1065 2535 -1055
rect 2600 -695 2650 -680
rect 2600 -1045 2610 -695
rect 2640 -1045 2650 -695
rect 2600 -1060 2650 -1045
rect 1720 -1280 1730 -1205
rect 1750 -1280 1760 -1205
rect 2605 -1135 2650 -1060
rect 2675 -685 2735 -620
rect 2675 -1055 2685 -685
rect 2725 -1055 2735 -685
rect 2675 -1065 2735 -1055
rect 2755 -685 2815 -620
rect 2755 -1055 2765 -685
rect 2805 -1055 2815 -685
rect 2755 -1065 2815 -1055
rect 2880 -695 2930 -680
rect 2880 -1045 2890 -695
rect 2920 -1045 2930 -695
rect 2880 -1060 2930 -1045
rect 2955 -685 3015 -620
rect 2955 -1055 2965 -685
rect 3005 -1055 3015 -685
rect 2885 -1135 2925 -1060
rect 2955 -1065 3015 -1055
rect 3040 -685 3100 -620
rect 3040 -1055 3050 -685
rect 3090 -1055 3100 -685
rect 3040 -1065 3100 -1055
rect 3165 -695 3215 -680
rect 3165 -1045 3175 -695
rect 3205 -1045 3215 -695
rect 3165 -1060 3215 -1045
rect 3240 -685 3300 -620
rect 3240 -1055 3250 -685
rect 3290 -1055 3300 -685
rect 3170 -1135 3210 -1060
rect 3240 -1065 3300 -1055
rect 3325 -685 3385 -620
rect 3325 -1055 3335 -685
rect 3375 -1055 3385 -685
rect 3325 -1065 3385 -1055
rect 3450 -695 3500 -680
rect 3450 -1045 3460 -695
rect 3490 -1045 3500 -695
rect 3450 -1060 3500 -1045
rect 3525 -685 3585 -620
rect 3525 -1055 3535 -685
rect 3575 -1055 3585 -685
rect 2605 -1145 2870 -1135
rect 2605 -1175 2790 -1145
rect 2860 -1175 2870 -1145
rect 2605 -1185 2870 -1175
rect 2885 -1145 3155 -1135
rect 2885 -1175 3075 -1145
rect 3145 -1175 3155 -1145
rect 2885 -1185 3155 -1175
rect 3170 -1145 3440 -1135
rect 3170 -1175 3360 -1145
rect 3430 -1175 3440 -1145
rect 3170 -1185 3440 -1175
rect 1720 -1285 1760 -1280
rect 2145 -1295 2195 -1265
rect 1435 -1320 1595 -1310
rect 1435 -1340 1540 -1320
rect 1585 -1340 1595 -1320
rect 1435 -1350 1595 -1340
rect 1885 -1360 1980 -1340
rect 1125 -1365 1420 -1360
rect 1610 -1365 1900 -1360
rect 1125 -1385 1900 -1365
rect 1965 -1385 1980 -1360
rect 2145 -1350 2155 -1295
rect 2185 -1340 2195 -1295
rect 2275 -1275 2580 -1265
rect 2275 -1300 2285 -1275
rect 2335 -1295 2530 -1275
rect 2570 -1295 2580 -1275
rect 2335 -1300 2580 -1295
rect 2275 -1305 2580 -1300
rect 2275 -1320 2325 -1305
rect 2520 -1340 2580 -1335
rect 2185 -1345 2580 -1340
rect 2185 -1350 2530 -1345
rect 2145 -1365 2530 -1350
rect 2570 -1365 2580 -1345
rect 2145 -1380 2580 -1365
rect 1125 -1400 1980 -1385
rect 2415 -1410 2585 -1395
rect 2415 -1415 2505 -1410
rect 1125 -1420 2505 -1415
rect 1125 -1445 1300 -1420
rect 1365 -1435 2505 -1420
rect 2570 -1435 2585 -1410
rect 1365 -1445 2585 -1435
rect 1125 -1455 2585 -1445
rect 1395 -1495 1475 -1480
rect 1395 -1750 1405 -1495
rect 1465 -1750 1475 -1495
rect 1395 -1835 1475 -1750
rect 1695 -1495 1775 -1480
rect 1695 -1750 1705 -1495
rect 1765 -1750 1775 -1495
rect 1695 -1835 1775 -1750
rect 1995 -1495 2075 -1480
rect 1995 -1750 2005 -1495
rect 2065 -1750 2075 -1495
rect 1995 -1835 2075 -1750
rect 2295 -1495 2375 -1480
rect 2295 -1750 2305 -1495
rect 2365 -1750 2375 -1495
rect 2295 -1835 2375 -1750
rect 2395 -1495 2475 -1480
rect 2605 -1485 2650 -1185
rect 2885 -1335 2925 -1185
rect 3170 -1265 3210 -1185
rect 2945 -1275 3210 -1265
rect 2945 -1295 2955 -1275
rect 2995 -1295 3210 -1275
rect 2945 -1305 3210 -1295
rect 2675 -1345 2925 -1335
rect 2675 -1365 2685 -1345
rect 2725 -1365 2925 -1345
rect 2675 -1375 2925 -1365
rect 2395 -1750 2405 -1495
rect 2465 -1750 2475 -1495
rect 2395 -1835 2475 -1750
rect 2600 -1500 2670 -1485
rect 2600 -1745 2610 -1500
rect 2660 -1745 2670 -1500
rect 2600 -1755 2670 -1745
rect 2754 -1495 2814 -1476
rect 2885 -1480 2925 -1375
rect 2754 -1645 2770 -1495
rect 2800 -1645 2814 -1495
rect 2754 -1835 2814 -1645
rect 2880 -1495 2930 -1480
rect 2880 -1645 2890 -1495
rect 2920 -1645 2930 -1495
rect 2880 -1660 2930 -1645
rect 2955 -1495 3015 -1475
rect 2955 -1645 2970 -1495
rect 3000 -1645 3015 -1495
rect 2955 -1835 3015 -1645
rect 3039 -1498 3099 -1475
rect 3170 -1480 3210 -1305
rect 3455 -1210 3495 -1060
rect 3525 -1065 3585 -1055
rect 3455 -1260 3620 -1210
rect 3039 -1648 3055 -1498
rect 3085 -1648 3099 -1498
rect 3039 -1835 3099 -1648
rect 3165 -1495 3215 -1480
rect 3165 -1645 3175 -1495
rect 3205 -1645 3215 -1495
rect 3165 -1660 3215 -1645
rect 3240 -1491 3300 -1475
rect 3240 -1641 3255 -1491
rect 3285 -1641 3300 -1491
rect 3240 -1835 3300 -1641
rect 3326 -1496 3386 -1475
rect 3455 -1480 3495 -1260
rect 3326 -1646 3339 -1496
rect 3369 -1646 3386 -1496
rect 3326 -1835 3386 -1646
rect 3450 -1495 3500 -1480
rect 3450 -1645 3460 -1495
rect 3490 -1645 3500 -1495
rect 3450 -1660 3500 -1645
rect 3525 -1493 3585 -1475
rect 3525 -1643 3541 -1493
rect 3571 -1643 3585 -1493
rect 3525 -1835 3585 -1643
rect 1125 -1895 3620 -1835
rect 1165 -2050 3580 -1895
rect 1005 -2070 3725 -2050
rect 1005 -2200 1050 -2070
rect 3695 -2200 3725 -2070
rect 1005 -2220 3725 -2200
<< via1 >>
rect 1255 -5 1305 40
rect 1355 -5 1405 40
rect 1455 -5 1505 40
rect 1555 -5 1605 40
rect 1655 -5 1705 40
rect 1755 -5 1805 40
rect 1855 -5 1905 40
rect 1955 -5 2005 40
rect 2055 -5 2105 40
rect 2155 -5 2205 40
rect 2255 -5 2305 40
rect 2355 -5 2405 40
rect 2455 -5 2505 40
rect 2555 -5 2605 40
rect 2655 -5 2705 40
rect 2755 -5 2805 40
rect 2855 -5 2905 40
rect 2955 -5 3005 40
rect 3055 -5 3105 40
rect 3155 -5 3205 40
rect 3255 -5 3305 40
rect 3355 -5 3405 40
rect 3455 -5 3505 40
rect 1255 -80 1305 -35
rect 1355 -80 1405 -35
rect 1455 -80 1505 -35
rect 1555 -80 1605 -35
rect 1655 -80 1705 -35
rect 1755 -80 1805 -35
rect 1855 -80 1905 -35
rect 1955 -80 2005 -35
rect 2055 -80 2105 -35
rect 2155 -80 2205 -35
rect 2255 -80 2305 -35
rect 2355 -80 2405 -35
rect 2455 -80 2505 -35
rect 2555 -80 2605 -35
rect 2655 -80 2705 -35
rect 2755 -80 2805 -35
rect 2855 -80 2905 -35
rect 2955 -80 3005 -35
rect 3055 -80 3105 -35
rect 3155 -80 3205 -35
rect 3255 -80 3305 -35
rect 3355 -80 3405 -35
rect 3455 -80 3505 -35
rect 1255 -155 1305 -110
rect 1355 -155 1405 -110
rect 1455 -155 1505 -110
rect 1555 -155 1605 -110
rect 1655 -155 1705 -110
rect 1755 -155 1805 -110
rect 1855 -155 1905 -110
rect 1955 -155 2005 -110
rect 2055 -155 2105 -110
rect 2155 -155 2205 -110
rect 2255 -155 2305 -110
rect 2355 -155 2405 -110
rect 2455 -155 2505 -110
rect 2555 -155 2605 -110
rect 2655 -155 2705 -110
rect 2755 -155 2805 -110
rect 2855 -155 2905 -110
rect 2955 -155 3005 -110
rect 3055 -155 3105 -110
rect 3155 -155 3205 -110
rect 3255 -155 3305 -110
rect 3355 -155 3405 -110
rect 3455 -155 3505 -110
rect 1050 -2200 3695 -2070
<< metal2 >>
rect 1200 40 3585 90
rect 1200 -5 1255 40
rect 1305 -5 1355 40
rect 1405 -5 1455 40
rect 1505 -5 1555 40
rect 1605 -5 1655 40
rect 1705 -5 1755 40
rect 1805 -5 1855 40
rect 1905 -5 1955 40
rect 2005 -5 2055 40
rect 2105 -5 2155 40
rect 2205 -5 2255 40
rect 2305 -5 2355 40
rect 2405 -5 2455 40
rect 2505 -5 2555 40
rect 2605 -5 2655 40
rect 2705 -5 2755 40
rect 2805 -5 2855 40
rect 2905 -5 2955 40
rect 3005 -5 3055 40
rect 3105 -5 3155 40
rect 3205 -5 3255 40
rect 3305 -5 3355 40
rect 3405 -5 3455 40
rect 3505 -5 3585 40
rect 1200 -35 3585 -5
rect 1200 -80 1255 -35
rect 1305 -80 1355 -35
rect 1405 -80 1455 -35
rect 1505 -80 1555 -35
rect 1605 -80 1655 -35
rect 1705 -80 1755 -35
rect 1805 -80 1855 -35
rect 1905 -80 1955 -35
rect 2005 -80 2055 -35
rect 2105 -80 2155 -35
rect 2205 -80 2255 -35
rect 2305 -80 2355 -35
rect 2405 -80 2455 -35
rect 2505 -80 2555 -35
rect 2605 -80 2655 -35
rect 2705 -80 2755 -35
rect 2805 -80 2855 -35
rect 2905 -80 2955 -35
rect 3005 -80 3055 -35
rect 3105 -80 3155 -35
rect 3205 -80 3255 -35
rect 3305 -80 3355 -35
rect 3405 -80 3455 -35
rect 3505 -80 3585 -35
rect 1200 -110 3585 -80
rect 1200 -155 1255 -110
rect 1305 -155 1355 -110
rect 1405 -155 1455 -110
rect 1505 -155 1555 -110
rect 1605 -155 1655 -110
rect 1705 -155 1755 -110
rect 1805 -155 1855 -110
rect 1905 -155 1955 -110
rect 2005 -155 2055 -110
rect 2105 -155 2155 -110
rect 2205 -155 2255 -110
rect 2305 -155 2355 -110
rect 2405 -155 2455 -110
rect 2505 -155 2555 -110
rect 2605 -155 2655 -110
rect 2705 -155 2755 -110
rect 2805 -155 2855 -110
rect 2905 -155 2955 -110
rect 3005 -155 3055 -110
rect 3105 -155 3155 -110
rect 3205 -155 3255 -110
rect 3305 -155 3355 -110
rect 3405 -155 3455 -110
rect 3505 -155 3585 -110
rect 1200 -190 3585 -155
rect 1005 -2070 3725 -2050
rect 1005 -2200 1050 -2070
rect 3695 -2200 3725 -2070
rect 1005 -2220 3725 -2200
<< via2 >>
rect 1255 -5 1305 40
rect 1355 -5 1405 40
rect 1455 -5 1505 40
rect 1555 -5 1605 40
rect 1655 -5 1705 40
rect 1755 -5 1805 40
rect 1855 -5 1905 40
rect 1955 -5 2005 40
rect 2055 -5 2105 40
rect 2155 -5 2205 40
rect 2255 -5 2305 40
rect 2355 -5 2405 40
rect 2455 -5 2505 40
rect 2555 -5 2605 40
rect 2655 -5 2705 40
rect 2755 -5 2805 40
rect 2855 -5 2905 40
rect 2955 -5 3005 40
rect 3055 -5 3105 40
rect 3155 -5 3205 40
rect 3255 -5 3305 40
rect 3355 -5 3405 40
rect 3455 -5 3505 40
rect 1255 -80 1305 -35
rect 1355 -80 1405 -35
rect 1455 -80 1505 -35
rect 1555 -80 1605 -35
rect 1655 -80 1705 -35
rect 1755 -80 1805 -35
rect 1855 -80 1905 -35
rect 1955 -80 2005 -35
rect 2055 -80 2105 -35
rect 2155 -80 2205 -35
rect 2255 -80 2305 -35
rect 2355 -80 2405 -35
rect 2455 -80 2505 -35
rect 2555 -80 2605 -35
rect 2655 -80 2705 -35
rect 2755 -80 2805 -35
rect 2855 -80 2905 -35
rect 2955 -80 3005 -35
rect 3055 -80 3105 -35
rect 3155 -80 3205 -35
rect 3255 -80 3305 -35
rect 3355 -80 3405 -35
rect 3455 -80 3505 -35
rect 1255 -155 1305 -110
rect 1355 -155 1405 -110
rect 1455 -155 1505 -110
rect 1555 -155 1605 -110
rect 1655 -155 1705 -110
rect 1755 -155 1805 -110
rect 1855 -155 1905 -110
rect 1955 -155 2005 -110
rect 2055 -155 2105 -110
rect 2155 -155 2205 -110
rect 2255 -155 2305 -110
rect 2355 -155 2405 -110
rect 2455 -155 2505 -110
rect 2555 -155 2605 -110
rect 2655 -155 2705 -110
rect 2755 -155 2805 -110
rect 2855 -155 2905 -110
rect 2955 -155 3005 -110
rect 3055 -155 3105 -110
rect 3155 -155 3205 -110
rect 3255 -155 3305 -110
rect 3355 -155 3405 -110
rect 3455 -155 3505 -110
rect 1050 -2200 3695 -2070
<< metal3 >>
rect 1200 40 3585 90
rect 1200 -5 1255 40
rect 1305 -5 1355 40
rect 1405 -5 1455 40
rect 1505 -5 1555 40
rect 1605 -5 1655 40
rect 1705 -5 1755 40
rect 1805 -5 1855 40
rect 1905 -5 1955 40
rect 2005 -5 2055 40
rect 2105 -5 2155 40
rect 2205 -5 2255 40
rect 2305 -5 2355 40
rect 2405 -5 2455 40
rect 2505 -5 2555 40
rect 2605 -5 2655 40
rect 2705 -5 2755 40
rect 2805 -5 2855 40
rect 2905 -5 2955 40
rect 3005 -5 3055 40
rect 3105 -5 3155 40
rect 3205 -5 3255 40
rect 3305 -5 3355 40
rect 3405 -5 3455 40
rect 3505 -5 3585 40
rect 1200 -35 3585 -5
rect 1200 -80 1255 -35
rect 1305 -80 1355 -35
rect 1405 -80 1455 -35
rect 1505 -80 1555 -35
rect 1605 -80 1655 -35
rect 1705 -80 1755 -35
rect 1805 -80 1855 -35
rect 1905 -80 1955 -35
rect 2005 -80 2055 -35
rect 2105 -80 2155 -35
rect 2205 -80 2255 -35
rect 2305 -80 2355 -35
rect 2405 -80 2455 -35
rect 2505 -80 2555 -35
rect 2605 -80 2655 -35
rect 2705 -80 2755 -35
rect 2805 -80 2855 -35
rect 2905 -80 2955 -35
rect 3005 -80 3055 -35
rect 3105 -80 3155 -35
rect 3205 -80 3255 -35
rect 3305 -80 3355 -35
rect 3405 -80 3455 -35
rect 3505 -80 3585 -35
rect 1200 -110 3585 -80
rect 1200 -155 1255 -110
rect 1305 -155 1355 -110
rect 1405 -155 1455 -110
rect 1505 -155 1555 -110
rect 1605 -155 1655 -110
rect 1705 -155 1755 -110
rect 1805 -155 1855 -110
rect 1905 -155 1955 -110
rect 2005 -155 2055 -110
rect 2105 -155 2155 -110
rect 2205 -155 2255 -110
rect 2305 -155 2355 -110
rect 2405 -155 2455 -110
rect 2505 -155 2555 -110
rect 2605 -155 2655 -110
rect 2705 -155 2755 -110
rect 2805 -155 2855 -110
rect 2905 -155 2955 -110
rect 3005 -155 3055 -110
rect 3105 -155 3155 -110
rect 3205 -155 3255 -110
rect 3305 -155 3355 -110
rect 3405 -155 3455 -110
rect 3505 -155 3585 -110
rect 1200 -190 3585 -155
rect 1005 -2070 3725 -2050
rect 1005 -2200 1050 -2070
rect 3695 -2200 3725 -2070
rect 1005 -2220 3725 -2200
<< via3 >>
rect 1050 -2200 3695 -2070
<< metal4 >>
rect 665 -495 4065 -190
rect 665 -1985 965 -495
rect 3765 -1985 4065 -495
rect 665 -2015 4065 -1985
rect 665 -2260 905 -2015
rect 965 -2050 3765 -2015
rect 950 -2070 3785 -2050
rect 950 -2200 1050 -2070
rect 3695 -2200 3785 -2070
rect 950 -2220 3785 -2200
rect 965 -2260 3765 -2220
rect 3815 -2260 4065 -2015
rect 665 -2290 4065 -2260
<< via4 >>
rect 1050 -2200 3695 -2070
<< metal5 >>
rect 665 -495 4065 -190
rect 665 -1985 965 -495
rect 3765 -1985 4065 -495
rect 665 -2070 4065 -1985
rect 665 -2200 1050 -2070
rect 3695 -2200 4065 -2070
rect 665 -2290 4065 -2200
<< labels >>
rlabel metal1 1125 -1254 1125 -1254 7 Vone
port 1 w
rlabel metal1 1125 -1147 1125 -1147 7 Vtwo
port 2 w
rlabel metal1 1125 -1381 1125 -1381 7 Ihyst
port 6 w
rlabel metal1 1125 -1436 1125 -1436 7 Ibias
port 3 w
rlabel metal1 3620 -1236 3620 -1236 3 OUT
port 7 e
rlabel metal1 1125 -1870 1125 -1870 7 VSS
port 4 w
rlabel metal1 1125 -590 1125 -590 7 VDD
port 5 w
<< end >>
