magic
tech sky130A
timestamp 1663665281
<< pwell >>
rect 169142 220939 169720 220950
rect 10383 219286 12006 220939
rect 32883 219286 34506 220939
rect 55383 219286 57006 220939
rect 77883 219286 79506 220939
rect 100383 219286 102006 220939
rect 122883 219286 124506 220939
rect 145383 219286 147006 220939
rect 167883 219286 169720 220939
rect 169142 219282 169720 219286
rect 189790 220115 192422 220956
rect 189790 220070 192265 220115
rect 192370 220070 192422 220115
rect 189790 219288 192422 220070
rect 189790 219285 191198 219288
rect 191820 219285 192422 219288
rect 208007 219036 219303 221128
rect 10383 196286 12006 197368
rect 32883 196286 34506 197368
rect 55383 196286 57006 197368
rect 77883 196286 79506 197368
rect 100383 196286 102006 197368
rect 122883 196286 124506 197368
rect 145383 196286 147006 197368
rect 167883 196286 169720 197368
rect 169142 196282 169720 196286
rect 189790 196288 192422 197368
rect 189790 196285 191198 196288
rect 191820 196285 192422 196288
rect 208007 196036 219303 197368
rect 10383 173286 12006 174368
rect 32883 173286 34506 174368
rect 55383 173286 57006 174368
rect 77883 173286 79506 174368
rect 100383 173286 102006 174368
rect 122883 173286 124506 174368
rect 145383 173286 147006 174368
rect 167883 173286 169720 174368
rect 169142 173282 169720 173286
rect 189790 173288 192422 174368
rect 189790 173285 191198 173288
rect 191820 173285 192422 173288
rect 208007 173036 219303 174368
rect 10383 150286 12006 151368
rect 32883 150286 34506 151368
rect 55383 150286 57006 151368
rect 77883 150286 79506 151368
rect 100383 150286 102006 151368
rect 122883 150286 124506 151368
rect 145383 150286 147006 151368
rect 167883 150286 169720 151368
rect 169142 150282 169720 150286
rect 189790 150288 192422 151368
rect 189790 150285 191198 150288
rect 191820 150285 192422 150288
rect 208007 150036 219303 151368
rect 10383 127286 12006 128368
rect 32883 127286 34506 128368
rect 55383 127286 57006 128368
rect 77883 127286 79506 128368
rect 100383 127286 102006 128368
rect 122883 127286 124506 128368
rect 145383 127286 147006 128368
rect 167883 127286 169720 128368
rect 169142 127282 169720 127286
rect 189790 127288 192422 128368
rect 189790 127285 191198 127288
rect 191820 127285 192422 127288
rect 208007 127036 219303 128368
rect 10383 104286 12006 105368
rect 32883 104286 34506 105368
rect 55383 104286 57006 105368
rect 77883 104286 79506 105368
rect 100383 104286 102006 105368
rect 122883 104286 124506 105368
rect 145383 104286 147006 105368
rect 167883 104286 169720 105368
rect 169142 104282 169720 104286
rect 189790 104288 192422 105368
rect 189790 104285 191198 104288
rect 191820 104285 192422 104288
rect 208007 104036 219303 105368
rect 10383 81286 12006 82368
rect 32883 81286 34506 82368
rect 55383 81286 57006 82368
rect 77883 81286 79506 82368
rect 100383 81286 102006 82368
rect 122883 81286 124506 82368
rect 145383 81286 147006 82368
rect 167883 81286 169720 82368
rect 169142 81282 169720 81286
rect 189790 81288 192422 82368
rect 189790 81285 191198 81288
rect 191820 81285 192422 81288
rect 208007 81036 219303 82368
rect 10383 58286 12006 59368
rect 32883 58286 34506 59368
rect 55383 58286 57006 59368
rect 77883 58286 79506 59368
rect 100383 58286 102006 59368
rect 122883 58286 124506 59368
rect 145383 58286 147006 59368
rect 167883 58286 169720 59368
rect 168091 58285 168458 58286
rect 169142 58282 169720 58286
rect 189790 58288 192422 59368
rect 189790 58285 191198 58288
rect 191820 58285 192422 58288
rect 208007 58036 219303 59368
rect 10383 35286 12006 36368
rect 32883 35286 34506 36368
rect 55383 35286 57006 36368
rect 77883 35286 79506 36368
rect 100383 35286 102006 36368
rect 122883 35286 124506 36368
rect 145383 35286 147006 36368
rect 167883 35286 169720 36368
rect 169142 35282 169720 35286
rect 189790 35288 192422 36368
rect 189790 35285 191198 35288
rect 191820 35285 192422 35288
rect 208007 35036 219303 36368
rect 9698 2236 12404 13659
rect 32365 2417 35071 13840
rect 54912 2236 57618 13659
rect 77519 2236 80225 13659
rect 99885 2116 102591 13539
rect 122552 2236 125258 13659
rect 144979 2357 147685 13780
rect 167525 2357 170231 13780
rect 189044 2336 192946 13566
rect 207545 2373 219474 13510
<< nmoslvt >>
rect 11166 220074 11181 220116
rect 33666 220074 33685 220116
rect 56166 220074 56191 220116
rect 78666 220074 78716 220116
rect 101166 220074 101266 220116
rect 123666 220074 123866 220116
rect 146166 220074 146566 220116
rect 168666 220074 169466 220116
rect 190166 220074 192166 220116
rect 208666 220074 218666 220116
rect 11166 197061 11181 197116
rect 33666 197061 33685 197116
rect 56166 197061 56191 197116
rect 78666 197061 78716 197116
rect 101166 197061 101266 197116
rect 123666 197061 123866 197116
rect 146166 197061 146566 197116
rect 168666 197061 169466 197116
rect 190166 197061 192166 197116
rect 208666 197061 218666 197116
rect 11166 174052 11181 174116
rect 33666 174052 33685 174116
rect 56166 174052 56191 174116
rect 78666 174052 78716 174116
rect 101166 174052 101266 174116
rect 123666 174052 123866 174116
rect 146166 174052 146566 174116
rect 168666 174052 169466 174116
rect 190166 174052 192166 174116
rect 208666 174052 218666 174116
rect 11166 151032 11181 151116
rect 33666 151032 33685 151116
rect 56166 151032 56191 151116
rect 78666 151032 78716 151116
rect 101166 151032 101266 151116
rect 123666 151032 123866 151116
rect 146166 151032 146566 151116
rect 168666 151032 169466 151116
rect 190166 151032 192166 151116
rect 208666 151032 218666 151116
rect 11166 128016 11181 128116
rect 33666 128016 33685 128116
rect 56166 128016 56191 128116
rect 78666 128016 78716 128116
rect 101166 128016 101266 128116
rect 123666 128016 123866 128116
rect 146166 128016 146566 128116
rect 168666 128016 169466 128116
rect 190166 128016 192166 128116
rect 208666 128016 218666 128116
rect 11166 104951 11181 105116
rect 33666 104951 33685 105116
rect 56166 104951 56191 105116
rect 78666 104951 78716 105116
rect 101166 104951 101266 105116
rect 123666 104951 123866 105116
rect 146166 104951 146566 105116
rect 168666 104951 169466 105116
rect 190166 104951 192166 105116
rect 208666 104951 218666 105116
rect 11166 81816 11181 82116
rect 33666 81816 33685 82116
rect 56166 81816 56191 82116
rect 78666 81816 78716 82116
rect 101166 81816 101266 82116
rect 123666 81816 123866 82116
rect 146166 81816 146566 82116
rect 168666 81816 169466 82116
rect 190166 81816 192166 82116
rect 208666 81816 218666 82116
rect 11166 58616 11181 59116
rect 33666 58616 33685 59116
rect 56166 58616 56191 59116
rect 78666 58616 78716 59116
rect 101166 58616 101266 59116
rect 123666 58616 123866 59116
rect 146166 58616 146566 59116
rect 168666 58616 169466 59116
rect 190166 58616 192166 59116
rect 208666 58616 218666 59116
rect 11166 35416 11181 36116
rect 33666 35416 33685 36116
rect 56166 35416 56191 36116
rect 78666 35416 78716 36116
rect 101166 35416 101266 36116
rect 123666 35416 123866 36116
rect 146166 35416 146566 36116
rect 168666 35416 169466 36116
rect 190166 35416 192166 36116
rect 208666 35416 218666 36116
rect 11166 3116 11181 13116
rect 33666 3116 33685 13116
rect 56166 3116 56191 13116
rect 78666 3116 78716 13116
rect 101166 3116 101266 13116
rect 123666 3116 123866 13116
rect 146166 3116 146566 13116
rect 168666 3116 169466 13116
rect 190166 3116 192166 13116
rect 208666 3116 218666 13116
<< ndiff >>
rect 11066 220103 11166 220116
rect 11066 220086 11078 220103
rect 11154 220086 11166 220103
rect 11066 220074 11166 220086
rect 11181 220103 11281 220116
rect 11181 220086 11193 220103
rect 11269 220086 11281 220103
rect 11181 220074 11281 220086
rect 33566 220103 33666 220116
rect 33566 220086 33578 220103
rect 33654 220086 33666 220103
rect 33566 220074 33666 220086
rect 33685 220103 33784 220116
rect 33685 220086 33696 220103
rect 33772 220086 33784 220103
rect 33685 220074 33784 220086
rect 56066 220103 56166 220116
rect 56066 220086 56078 220103
rect 56154 220086 56166 220103
rect 56066 220074 56166 220086
rect 56191 220103 56291 220116
rect 56191 220086 56203 220103
rect 56279 220086 56291 220103
rect 56191 220074 56291 220086
rect 78566 220103 78666 220116
rect 78566 220086 78578 220103
rect 78654 220086 78666 220103
rect 78566 220074 78666 220086
rect 78716 220103 78816 220116
rect 78716 220086 78728 220103
rect 78804 220086 78816 220103
rect 78716 220074 78816 220086
rect 101066 220103 101166 220116
rect 101066 220086 101078 220103
rect 101154 220086 101166 220103
rect 101066 220074 101166 220086
rect 101266 220103 101366 220116
rect 101266 220086 101278 220103
rect 101354 220086 101366 220103
rect 101266 220074 101366 220086
rect 123566 220103 123666 220116
rect 123566 220086 123578 220103
rect 123654 220086 123666 220103
rect 123566 220074 123666 220086
rect 123866 220103 123966 220116
rect 123866 220086 123878 220103
rect 123954 220086 123966 220103
rect 123866 220074 123966 220086
rect 146066 220103 146166 220116
rect 146066 220086 146078 220103
rect 146154 220086 146166 220103
rect 146066 220074 146166 220086
rect 146566 220103 146666 220116
rect 146566 220086 146578 220103
rect 146654 220086 146666 220103
rect 146566 220074 146666 220086
rect 168566 220103 168666 220116
rect 168566 220086 168578 220103
rect 168654 220086 168666 220103
rect 168566 220074 168666 220086
rect 169466 220103 169566 220116
rect 169466 220086 169478 220103
rect 169554 220086 169566 220103
rect 169466 220074 169566 220086
rect 190066 220103 190166 220116
rect 190066 220086 190078 220103
rect 190154 220086 190166 220103
rect 190066 220074 190166 220086
rect 192166 220103 192266 220116
rect 192166 220086 192178 220103
rect 192254 220086 192266 220103
rect 192166 220074 192266 220086
rect 208566 220103 208666 220116
rect 208566 220086 208578 220103
rect 208654 220086 208666 220103
rect 208566 220074 208666 220086
rect 218666 220103 218766 220116
rect 218666 220086 218678 220103
rect 218754 220086 218766 220103
rect 218666 220074 218766 220086
rect 11066 197103 11166 197116
rect 11066 197073 11078 197103
rect 11154 197073 11166 197103
rect 11066 197061 11166 197073
rect 11181 197103 11281 197116
rect 11181 197073 11193 197103
rect 11269 197073 11281 197103
rect 11181 197061 11281 197073
rect 33566 197103 33666 197116
rect 33566 197073 33578 197103
rect 33654 197073 33666 197103
rect 33566 197061 33666 197073
rect 33685 197103 33784 197116
rect 33685 197073 33696 197103
rect 33772 197073 33784 197103
rect 33685 197061 33784 197073
rect 56066 197103 56166 197116
rect 56066 197073 56078 197103
rect 56154 197073 56166 197103
rect 56066 197061 56166 197073
rect 56191 197103 56291 197116
rect 56191 197073 56203 197103
rect 56279 197073 56291 197103
rect 56191 197061 56291 197073
rect 78566 197103 78666 197116
rect 78566 197073 78578 197103
rect 78654 197073 78666 197103
rect 78566 197061 78666 197073
rect 78716 197103 78816 197116
rect 78716 197073 78728 197103
rect 78804 197073 78816 197103
rect 78716 197061 78816 197073
rect 101066 197103 101166 197116
rect 101066 197073 101078 197103
rect 101154 197073 101166 197103
rect 101066 197061 101166 197073
rect 101266 197103 101366 197116
rect 101266 197073 101278 197103
rect 101354 197073 101366 197103
rect 101266 197061 101366 197073
rect 123566 197103 123666 197116
rect 123566 197073 123578 197103
rect 123654 197073 123666 197103
rect 123566 197061 123666 197073
rect 123866 197103 123966 197116
rect 123866 197073 123878 197103
rect 123954 197073 123966 197103
rect 123866 197061 123966 197073
rect 146066 197103 146166 197116
rect 146066 197073 146078 197103
rect 146154 197073 146166 197103
rect 146066 197061 146166 197073
rect 146566 197103 146666 197116
rect 146566 197073 146578 197103
rect 146654 197073 146666 197103
rect 146566 197061 146666 197073
rect 168566 197103 168666 197116
rect 168566 197073 168578 197103
rect 168654 197073 168666 197103
rect 168566 197061 168666 197073
rect 169466 197103 169566 197116
rect 169466 197073 169478 197103
rect 169554 197073 169566 197103
rect 169466 197061 169566 197073
rect 190066 197103 190166 197116
rect 190066 197073 190078 197103
rect 190154 197073 190166 197103
rect 190066 197061 190166 197073
rect 192166 197103 192266 197116
rect 192166 197073 192178 197103
rect 192254 197073 192266 197103
rect 192166 197061 192266 197073
rect 208566 197103 208666 197116
rect 208566 197073 208578 197103
rect 208654 197073 208666 197103
rect 208566 197061 208666 197073
rect 218666 197103 218766 197116
rect 218666 197073 218678 197103
rect 218754 197073 218766 197103
rect 218666 197061 218766 197073
rect 11066 174103 11166 174116
rect 11066 174064 11078 174103
rect 11154 174064 11166 174103
rect 11066 174052 11166 174064
rect 11181 174103 11281 174116
rect 11181 174064 11193 174103
rect 11269 174064 11281 174103
rect 11181 174052 11281 174064
rect 33566 174103 33666 174116
rect 33566 174064 33578 174103
rect 33654 174064 33666 174103
rect 33566 174052 33666 174064
rect 33685 174103 33784 174116
rect 33685 174064 33696 174103
rect 33772 174064 33784 174103
rect 33685 174052 33784 174064
rect 56066 174103 56166 174116
rect 56066 174064 56078 174103
rect 56154 174064 56166 174103
rect 56066 174052 56166 174064
rect 56191 174103 56291 174116
rect 56191 174064 56203 174103
rect 56279 174064 56291 174103
rect 56191 174052 56291 174064
rect 78566 174103 78666 174116
rect 78566 174064 78578 174103
rect 78654 174064 78666 174103
rect 78566 174052 78666 174064
rect 78716 174103 78816 174116
rect 78716 174064 78728 174103
rect 78804 174064 78816 174103
rect 78716 174052 78816 174064
rect 101066 174103 101166 174116
rect 101066 174064 101078 174103
rect 101154 174064 101166 174103
rect 101066 174052 101166 174064
rect 101266 174103 101366 174116
rect 101266 174064 101278 174103
rect 101354 174064 101366 174103
rect 101266 174052 101366 174064
rect 123566 174103 123666 174116
rect 123566 174064 123578 174103
rect 123654 174064 123666 174103
rect 123566 174052 123666 174064
rect 123866 174103 123966 174116
rect 123866 174064 123878 174103
rect 123954 174064 123966 174103
rect 123866 174052 123966 174064
rect 146066 174103 146166 174116
rect 146066 174064 146078 174103
rect 146154 174064 146166 174103
rect 146066 174052 146166 174064
rect 146566 174103 146666 174116
rect 146566 174064 146578 174103
rect 146654 174064 146666 174103
rect 146566 174052 146666 174064
rect 168566 174103 168666 174116
rect 168566 174064 168578 174103
rect 168654 174064 168666 174103
rect 168566 174052 168666 174064
rect 169466 174103 169566 174116
rect 169466 174064 169478 174103
rect 169554 174064 169566 174103
rect 169466 174052 169566 174064
rect 190066 174103 190166 174116
rect 190066 174064 190078 174103
rect 190154 174064 190166 174103
rect 190066 174052 190166 174064
rect 192166 174103 192266 174116
rect 192166 174064 192178 174103
rect 192254 174064 192266 174103
rect 192166 174052 192266 174064
rect 208566 174103 208666 174116
rect 208566 174064 208578 174103
rect 208654 174064 208666 174103
rect 208566 174052 208666 174064
rect 218666 174103 218766 174116
rect 218666 174064 218678 174103
rect 218754 174064 218766 174103
rect 218666 174052 218766 174064
rect 11066 151103 11166 151116
rect 11066 151044 11078 151103
rect 11154 151044 11166 151103
rect 11066 151032 11166 151044
rect 11181 151103 11281 151116
rect 11181 151044 11193 151103
rect 11269 151044 11281 151103
rect 11181 151032 11281 151044
rect 33566 151103 33666 151116
rect 33566 151044 33578 151103
rect 33654 151044 33666 151103
rect 33566 151032 33666 151044
rect 33685 151103 33784 151116
rect 33685 151044 33696 151103
rect 33772 151044 33784 151103
rect 33685 151032 33784 151044
rect 56066 151103 56166 151116
rect 56066 151044 56078 151103
rect 56154 151044 56166 151103
rect 56066 151032 56166 151044
rect 56191 151103 56291 151116
rect 56191 151044 56203 151103
rect 56279 151044 56291 151103
rect 56191 151032 56291 151044
rect 78566 151103 78666 151116
rect 78566 151044 78578 151103
rect 78654 151044 78666 151103
rect 78566 151032 78666 151044
rect 78716 151103 78816 151116
rect 78716 151044 78728 151103
rect 78804 151044 78816 151103
rect 78716 151032 78816 151044
rect 101066 151103 101166 151116
rect 101066 151044 101078 151103
rect 101154 151044 101166 151103
rect 101066 151032 101166 151044
rect 101266 151103 101366 151116
rect 101266 151044 101278 151103
rect 101354 151044 101366 151103
rect 101266 151032 101366 151044
rect 123566 151103 123666 151116
rect 123566 151044 123578 151103
rect 123654 151044 123666 151103
rect 123566 151032 123666 151044
rect 123866 151103 123966 151116
rect 123866 151044 123878 151103
rect 123954 151044 123966 151103
rect 123866 151032 123966 151044
rect 146066 151103 146166 151116
rect 146066 151044 146078 151103
rect 146154 151044 146166 151103
rect 146066 151032 146166 151044
rect 146566 151103 146666 151116
rect 146566 151044 146578 151103
rect 146654 151044 146666 151103
rect 146566 151032 146666 151044
rect 168566 151103 168666 151116
rect 168566 151044 168578 151103
rect 168654 151044 168666 151103
rect 168566 151032 168666 151044
rect 169466 151103 169566 151116
rect 169466 151044 169478 151103
rect 169554 151044 169566 151103
rect 169466 151032 169566 151044
rect 190066 151103 190166 151116
rect 190066 151044 190078 151103
rect 190154 151044 190166 151103
rect 190066 151032 190166 151044
rect 192166 151103 192266 151116
rect 192166 151044 192178 151103
rect 192254 151044 192266 151103
rect 192166 151032 192266 151044
rect 208566 151103 208666 151116
rect 208566 151044 208578 151103
rect 208654 151044 208666 151103
rect 208566 151032 208666 151044
rect 218666 151103 218766 151116
rect 218666 151044 218678 151103
rect 218754 151044 218766 151103
rect 218666 151032 218766 151044
rect 11066 128103 11166 128116
rect 11066 128028 11078 128103
rect 11154 128028 11166 128103
rect 11066 128016 11166 128028
rect 11181 128103 11281 128116
rect 11181 128028 11193 128103
rect 11269 128028 11281 128103
rect 11181 128016 11281 128028
rect 33566 128103 33666 128116
rect 33566 128028 33578 128103
rect 33654 128028 33666 128103
rect 33566 128016 33666 128028
rect 33685 128103 33784 128116
rect 33685 128028 33696 128103
rect 33772 128028 33784 128103
rect 33685 128016 33784 128028
rect 56066 128103 56166 128116
rect 56066 128028 56078 128103
rect 56154 128028 56166 128103
rect 56066 128016 56166 128028
rect 56191 128103 56291 128116
rect 56191 128028 56203 128103
rect 56279 128028 56291 128103
rect 56191 128016 56291 128028
rect 78566 128103 78666 128116
rect 78566 128028 78578 128103
rect 78654 128028 78666 128103
rect 78566 128016 78666 128028
rect 78716 128103 78816 128116
rect 78716 128028 78728 128103
rect 78804 128028 78816 128103
rect 78716 128016 78816 128028
rect 101066 128103 101166 128116
rect 101066 128028 101078 128103
rect 101154 128028 101166 128103
rect 101066 128016 101166 128028
rect 101266 128103 101366 128116
rect 101266 128028 101278 128103
rect 101354 128028 101366 128103
rect 101266 128016 101366 128028
rect 123566 128103 123666 128116
rect 123566 128028 123578 128103
rect 123654 128028 123666 128103
rect 123566 128016 123666 128028
rect 123866 128103 123966 128116
rect 123866 128028 123878 128103
rect 123954 128028 123966 128103
rect 123866 128016 123966 128028
rect 146066 128103 146166 128116
rect 146066 128028 146078 128103
rect 146154 128028 146166 128103
rect 146066 128016 146166 128028
rect 146566 128103 146666 128116
rect 146566 128028 146578 128103
rect 146654 128028 146666 128103
rect 146566 128016 146666 128028
rect 168566 128103 168666 128116
rect 168566 128028 168578 128103
rect 168654 128028 168666 128103
rect 168566 128016 168666 128028
rect 169466 128103 169566 128116
rect 169466 128028 169478 128103
rect 169554 128028 169566 128103
rect 169466 128016 169566 128028
rect 190066 128103 190166 128116
rect 190066 128028 190078 128103
rect 190154 128028 190166 128103
rect 190066 128016 190166 128028
rect 192166 128103 192266 128116
rect 192166 128028 192178 128103
rect 192254 128028 192266 128103
rect 192166 128016 192266 128028
rect 208566 128103 208666 128116
rect 208566 128028 208578 128103
rect 208654 128028 208666 128103
rect 208566 128016 208666 128028
rect 218666 128103 218766 128116
rect 218666 128028 218678 128103
rect 218754 128028 218766 128103
rect 218666 128016 218766 128028
rect 11066 105103 11166 105116
rect 11066 104963 11078 105103
rect 11154 104963 11166 105103
rect 11066 104951 11166 104963
rect 11181 105103 11281 105116
rect 11181 104963 11193 105103
rect 11269 104963 11281 105103
rect 11181 104951 11281 104963
rect 33566 105103 33666 105116
rect 33566 104963 33578 105103
rect 33654 104963 33666 105103
rect 33566 104951 33666 104963
rect 33685 105103 33784 105116
rect 33685 104963 33696 105103
rect 33772 104963 33784 105103
rect 33685 104951 33784 104963
rect 56066 105103 56166 105116
rect 56066 104963 56078 105103
rect 56154 104963 56166 105103
rect 56066 104951 56166 104963
rect 56191 105103 56291 105116
rect 56191 104963 56203 105103
rect 56279 104963 56291 105103
rect 56191 104951 56291 104963
rect 78566 105103 78666 105116
rect 78566 104963 78578 105103
rect 78654 104963 78666 105103
rect 78566 104951 78666 104963
rect 78716 105103 78816 105116
rect 78716 104963 78728 105103
rect 78804 104963 78816 105103
rect 78716 104951 78816 104963
rect 101066 105103 101166 105116
rect 101066 104963 101078 105103
rect 101154 104963 101166 105103
rect 101066 104951 101166 104963
rect 101266 105103 101366 105116
rect 101266 104963 101278 105103
rect 101354 104963 101366 105103
rect 101266 104951 101366 104963
rect 123566 105103 123666 105116
rect 123566 104963 123578 105103
rect 123654 104963 123666 105103
rect 123566 104951 123666 104963
rect 123866 105103 123966 105116
rect 123866 104963 123878 105103
rect 123954 104963 123966 105103
rect 123866 104951 123966 104963
rect 146066 105103 146166 105116
rect 146066 104963 146078 105103
rect 146154 104963 146166 105103
rect 146066 104951 146166 104963
rect 146566 105103 146666 105116
rect 146566 104963 146578 105103
rect 146654 104963 146666 105103
rect 146566 104951 146666 104963
rect 168566 105103 168666 105116
rect 168566 104963 168578 105103
rect 168654 104963 168666 105103
rect 168566 104951 168666 104963
rect 169466 105103 169566 105116
rect 169466 104963 169478 105103
rect 169554 104963 169566 105103
rect 169466 104951 169566 104963
rect 190066 105103 190166 105116
rect 190066 104963 190078 105103
rect 190154 104963 190166 105103
rect 190066 104951 190166 104963
rect 192166 105103 192266 105116
rect 192166 104963 192178 105103
rect 192254 104963 192266 105103
rect 192166 104951 192266 104963
rect 208566 105103 208666 105116
rect 208566 104963 208578 105103
rect 208654 104963 208666 105103
rect 208566 104951 208666 104963
rect 218666 105103 218766 105116
rect 218666 104963 218678 105103
rect 218754 104963 218766 105103
rect 218666 104951 218766 104963
rect 11066 82103 11166 82116
rect 11066 81828 11078 82103
rect 11154 81828 11166 82103
rect 11066 81816 11166 81828
rect 11181 82103 11281 82116
rect 11181 81828 11193 82103
rect 11269 81828 11281 82103
rect 11181 81816 11281 81828
rect 33566 82103 33666 82116
rect 33566 81828 33578 82103
rect 33654 81828 33666 82103
rect 33566 81816 33666 81828
rect 33685 82103 33784 82116
rect 33685 81828 33696 82103
rect 33772 81828 33784 82103
rect 33685 81816 33784 81828
rect 56066 82103 56166 82116
rect 56066 81828 56078 82103
rect 56154 81828 56166 82103
rect 56066 81816 56166 81828
rect 56191 82103 56291 82116
rect 56191 81828 56203 82103
rect 56279 81828 56291 82103
rect 56191 81816 56291 81828
rect 78566 82103 78666 82116
rect 78566 81828 78578 82103
rect 78654 81828 78666 82103
rect 78566 81816 78666 81828
rect 78716 82103 78816 82116
rect 78716 81828 78728 82103
rect 78804 81828 78816 82103
rect 78716 81816 78816 81828
rect 101066 82103 101166 82116
rect 101066 81828 101078 82103
rect 101154 81828 101166 82103
rect 101066 81816 101166 81828
rect 101266 82103 101366 82116
rect 101266 81828 101278 82103
rect 101354 81828 101366 82103
rect 101266 81816 101366 81828
rect 123566 82103 123666 82116
rect 123566 81828 123578 82103
rect 123654 81828 123666 82103
rect 123566 81816 123666 81828
rect 123866 82103 123966 82116
rect 123866 81828 123878 82103
rect 123954 81828 123966 82103
rect 123866 81816 123966 81828
rect 146066 82103 146166 82116
rect 146066 81828 146078 82103
rect 146154 81828 146166 82103
rect 146066 81816 146166 81828
rect 146566 82103 146666 82116
rect 146566 81828 146578 82103
rect 146654 81828 146666 82103
rect 146566 81816 146666 81828
rect 168566 82103 168666 82116
rect 168566 81828 168578 82103
rect 168654 81828 168666 82103
rect 168566 81816 168666 81828
rect 169466 82103 169566 82116
rect 169466 81828 169478 82103
rect 169554 81828 169566 82103
rect 169466 81816 169566 81828
rect 190066 82103 190166 82116
rect 190066 81828 190078 82103
rect 190154 81828 190166 82103
rect 190066 81816 190166 81828
rect 192166 82103 192266 82116
rect 192166 81828 192178 82103
rect 192254 81828 192266 82103
rect 192166 81816 192266 81828
rect 208566 82103 208666 82116
rect 208566 81828 208578 82103
rect 208654 81828 208666 82103
rect 208566 81816 208666 81828
rect 218666 82103 218766 82116
rect 218666 81828 218678 82103
rect 218754 81828 218766 82103
rect 218666 81816 218766 81828
rect 11066 59103 11166 59116
rect 11066 58628 11078 59103
rect 11154 58628 11166 59103
rect 11066 58616 11166 58628
rect 11181 59103 11281 59116
rect 11181 58628 11193 59103
rect 11269 58946 11281 59103
rect 11275 58633 11281 58946
rect 11269 58628 11281 58633
rect 11181 58616 11281 58628
rect 33566 59103 33666 59116
rect 33566 58628 33578 59103
rect 33654 58628 33666 59103
rect 33566 58616 33666 58628
rect 33685 59103 33784 59116
rect 33685 58628 33696 59103
rect 33772 58628 33784 59103
rect 33685 58616 33784 58628
rect 56066 59103 56166 59116
rect 56066 58628 56078 59103
rect 56154 58628 56166 59103
rect 56066 58616 56166 58628
rect 56191 59103 56291 59116
rect 56191 58628 56203 59103
rect 56279 58628 56291 59103
rect 56191 58616 56291 58628
rect 78566 59103 78666 59116
rect 78566 58628 78578 59103
rect 78654 58628 78666 59103
rect 78566 58616 78666 58628
rect 78716 59103 78816 59116
rect 78716 58628 78728 59103
rect 78804 58628 78816 59103
rect 78716 58616 78816 58628
rect 101066 59103 101166 59116
rect 101066 58628 101078 59103
rect 101154 58628 101166 59103
rect 101066 58616 101166 58628
rect 101266 59103 101366 59116
rect 101266 58628 101278 59103
rect 101354 58628 101366 59103
rect 101266 58616 101366 58628
rect 123566 59103 123666 59116
rect 123566 58628 123578 59103
rect 123654 58628 123666 59103
rect 123566 58616 123666 58628
rect 123866 59103 123966 59116
rect 123866 58628 123878 59103
rect 123954 58628 123966 59103
rect 146066 59103 146166 59116
rect 123866 58616 123966 58628
rect 146066 58628 146078 59103
rect 146154 58628 146166 59103
rect 146066 58616 146166 58628
rect 146566 59103 146666 59116
rect 146566 58628 146578 59103
rect 146654 58628 146666 59103
rect 146566 58616 146666 58628
rect 168566 59103 168666 59116
rect 168566 58628 168578 59103
rect 168654 58628 168666 59103
rect 168566 58616 168666 58628
rect 169466 59103 169566 59116
rect 169466 58628 169478 59103
rect 169554 58628 169566 59103
rect 169466 58616 169566 58628
rect 190066 59103 190166 59116
rect 190066 58628 190078 59103
rect 190154 58628 190166 59103
rect 190066 58616 190166 58628
rect 192166 59103 192266 59116
rect 192166 58628 192178 59103
rect 192254 58628 192266 59103
rect 192166 58616 192266 58628
rect 208566 59103 208666 59116
rect 208566 58628 208578 59103
rect 208654 58628 208666 59103
rect 208566 58616 208666 58628
rect 218666 59103 218766 59116
rect 218666 58628 218678 59103
rect 218754 58628 218766 59103
rect 218666 58616 218766 58628
rect 11066 36103 11166 36116
rect 11066 35428 11078 36103
rect 11154 35428 11166 36103
rect 11066 35416 11166 35428
rect 11181 36103 11281 36116
rect 11181 35428 11193 36103
rect 11269 35428 11281 36103
rect 11181 35416 11281 35428
rect 33566 36103 33666 36116
rect 33566 35428 33578 36103
rect 33654 35428 33666 36103
rect 33566 35416 33666 35428
rect 33685 36103 33784 36116
rect 33685 35428 33696 36103
rect 33772 35428 33784 36103
rect 33685 35416 33784 35428
rect 56066 36103 56166 36116
rect 56066 35428 56078 36103
rect 56154 35428 56166 36103
rect 56066 35416 56166 35428
rect 56191 36103 56291 36116
rect 56191 35428 56203 36103
rect 56279 35428 56291 36103
rect 56191 35416 56291 35428
rect 78566 36103 78666 36116
rect 78566 35428 78578 36103
rect 78654 35428 78666 36103
rect 78566 35416 78666 35428
rect 78716 36103 78816 36116
rect 78716 35428 78728 36103
rect 78804 35428 78816 36103
rect 78716 35416 78816 35428
rect 101066 36103 101166 36116
rect 101066 35428 101078 36103
rect 101154 35428 101166 36103
rect 101066 35416 101166 35428
rect 101266 36103 101366 36116
rect 101266 35428 101278 36103
rect 101354 35428 101366 36103
rect 101266 35416 101366 35428
rect 123566 36103 123666 36116
rect 123566 35428 123578 36103
rect 123654 35428 123666 36103
rect 123566 35416 123666 35428
rect 123866 36103 123966 36116
rect 123866 35428 123878 36103
rect 123954 35428 123966 36103
rect 123866 35416 123966 35428
rect 146066 36103 146166 36116
rect 146066 35428 146078 36103
rect 146154 35428 146166 36103
rect 146066 35416 146166 35428
rect 146566 36103 146666 36116
rect 146566 35428 146578 36103
rect 146654 35428 146666 36103
rect 146566 35416 146666 35428
rect 168566 36103 168666 36116
rect 168566 35428 168578 36103
rect 168654 35428 168666 36103
rect 168566 35416 168666 35428
rect 169466 36103 169566 36116
rect 169466 35428 169478 36103
rect 169554 35428 169566 36103
rect 169466 35416 169566 35428
rect 190066 36103 190166 36116
rect 190066 35428 190078 36103
rect 190154 35428 190166 36103
rect 190066 35416 190166 35428
rect 192166 36103 192266 36116
rect 192166 35428 192178 36103
rect 192254 35428 192266 36103
rect 192166 35416 192266 35428
rect 208566 36103 208666 36116
rect 208566 35428 208578 36103
rect 208654 35428 208666 36103
rect 208566 35416 208666 35428
rect 218666 36103 218766 36116
rect 218666 35428 218678 36103
rect 218754 35428 218766 36103
rect 218666 35416 218766 35428
rect 11066 13103 11166 13116
rect 11066 3128 11078 13103
rect 11154 3128 11166 13103
rect 11066 3116 11166 3128
rect 11181 13103 11281 13116
rect 11181 3128 11193 13103
rect 11269 3128 11281 13103
rect 11181 3116 11281 3128
rect 33566 13103 33666 13116
rect 33566 3128 33578 13103
rect 33654 3128 33666 13103
rect 33566 3116 33666 3128
rect 33685 13103 33784 13116
rect 33685 3128 33696 13103
rect 33772 3128 33784 13103
rect 33685 3116 33784 3128
rect 56066 13103 56166 13116
rect 56066 3128 56078 13103
rect 56154 3128 56166 13103
rect 56066 3116 56166 3128
rect 56191 13103 56291 13116
rect 56191 3128 56203 13103
rect 56279 3128 56291 13103
rect 56191 3116 56291 3128
rect 78566 13103 78666 13116
rect 78566 3128 78578 13103
rect 78654 3128 78666 13103
rect 78566 3116 78666 3128
rect 78716 13103 78816 13116
rect 78716 3128 78728 13103
rect 78804 3128 78816 13103
rect 78716 3116 78816 3128
rect 101066 13103 101166 13116
rect 101066 3128 101078 13103
rect 101154 3128 101166 13103
rect 101066 3116 101166 3128
rect 101266 13103 101366 13116
rect 101266 3128 101278 13103
rect 101354 3128 101366 13103
rect 101266 3116 101366 3128
rect 123566 13103 123666 13116
rect 123566 3128 123578 13103
rect 123654 3128 123666 13103
rect 123566 3116 123666 3128
rect 123866 13103 123966 13116
rect 123866 3128 123878 13103
rect 123954 3128 123966 13103
rect 123866 3116 123966 3128
rect 146066 13103 146166 13116
rect 146066 3128 146078 13103
rect 146154 3128 146166 13103
rect 146066 3116 146166 3128
rect 146566 13103 146666 13116
rect 146566 3128 146578 13103
rect 146654 3128 146666 13103
rect 146566 3116 146666 3128
rect 168566 13103 168666 13116
rect 168566 3128 168578 13103
rect 168654 3128 168666 13103
rect 168566 3116 168666 3128
rect 169466 13103 169566 13116
rect 169466 3128 169478 13103
rect 169554 3128 169566 13103
rect 169466 3116 169566 3128
rect 190066 13103 190166 13116
rect 190066 3128 190078 13103
rect 190154 3128 190166 13103
rect 190066 3116 190166 3128
rect 192166 13103 192266 13116
rect 192166 3128 192178 13103
rect 192254 3128 192266 13103
rect 192166 3116 192266 3128
rect 208566 13103 208666 13116
rect 208566 3128 208578 13103
rect 208654 3128 208666 13103
rect 208566 3116 208666 3128
rect 218666 13103 218766 13116
rect 218666 3128 218678 13103
rect 218754 3128 218766 13103
rect 218666 3116 218766 3128
<< ndiffc >>
rect 11078 220086 11154 220103
rect 11193 220086 11269 220103
rect 33578 220086 33654 220103
rect 33696 220086 33772 220103
rect 56078 220086 56154 220103
rect 56203 220086 56279 220103
rect 78578 220086 78654 220103
rect 78728 220086 78804 220103
rect 101078 220086 101154 220103
rect 101278 220086 101354 220103
rect 123578 220086 123654 220103
rect 123878 220086 123954 220103
rect 146078 220086 146154 220103
rect 146578 220086 146654 220103
rect 168578 220086 168654 220103
rect 169478 220086 169554 220103
rect 190078 220086 190154 220103
rect 192178 220086 192254 220103
rect 208578 220086 208654 220103
rect 218678 220086 218754 220103
rect 11078 197073 11154 197103
rect 11193 197073 11269 197103
rect 33578 197073 33654 197103
rect 33696 197073 33772 197103
rect 56078 197073 56154 197103
rect 56203 197073 56279 197103
rect 78578 197073 78654 197103
rect 78728 197073 78804 197103
rect 101078 197073 101154 197103
rect 101278 197073 101354 197103
rect 123578 197073 123654 197103
rect 123878 197073 123954 197103
rect 146078 197073 146154 197103
rect 146578 197073 146654 197103
rect 168578 197073 168654 197103
rect 169478 197073 169554 197103
rect 190078 197073 190154 197103
rect 192178 197073 192254 197103
rect 208578 197073 208654 197103
rect 218678 197073 218754 197103
rect 11078 174064 11154 174103
rect 11193 174064 11269 174103
rect 33578 174064 33654 174103
rect 33696 174064 33772 174103
rect 56078 174064 56154 174103
rect 56203 174064 56279 174103
rect 78578 174064 78654 174103
rect 78728 174064 78804 174103
rect 101078 174064 101154 174103
rect 101278 174064 101354 174103
rect 123578 174064 123654 174103
rect 123878 174064 123954 174103
rect 146078 174064 146154 174103
rect 146578 174064 146654 174103
rect 168578 174064 168654 174103
rect 169478 174064 169554 174103
rect 190078 174064 190154 174103
rect 192178 174064 192254 174103
rect 208578 174064 208654 174103
rect 218678 174064 218754 174103
rect 11078 151044 11154 151103
rect 11193 151044 11269 151103
rect 33578 151044 33654 151103
rect 33696 151044 33772 151103
rect 56078 151044 56154 151103
rect 56203 151044 56279 151103
rect 78578 151044 78654 151103
rect 78728 151044 78804 151103
rect 101078 151044 101154 151103
rect 101278 151044 101354 151103
rect 123578 151044 123654 151103
rect 123878 151044 123954 151103
rect 146078 151044 146154 151103
rect 146578 151044 146654 151103
rect 168578 151044 168654 151103
rect 169478 151044 169554 151103
rect 190078 151044 190154 151103
rect 192178 151044 192254 151103
rect 208578 151044 208654 151103
rect 218678 151044 218754 151103
rect 11078 128028 11154 128103
rect 11193 128028 11269 128103
rect 33578 128028 33654 128103
rect 33696 128028 33772 128103
rect 56078 128028 56154 128103
rect 56203 128028 56279 128103
rect 78578 128028 78654 128103
rect 78728 128028 78804 128103
rect 101078 128028 101154 128103
rect 101278 128028 101354 128103
rect 123578 128028 123654 128103
rect 123878 128028 123954 128103
rect 146078 128028 146154 128103
rect 146578 128028 146654 128103
rect 168578 128028 168654 128103
rect 169478 128028 169554 128103
rect 190078 128028 190154 128103
rect 192178 128028 192254 128103
rect 208578 128028 208654 128103
rect 218678 128028 218754 128103
rect 11078 104963 11154 105103
rect 11193 104963 11269 105103
rect 33578 104963 33654 105103
rect 33696 104963 33772 105103
rect 56078 104963 56154 105103
rect 56203 104963 56279 105103
rect 78578 104963 78654 105103
rect 78728 104963 78804 105103
rect 101078 104963 101154 105103
rect 101278 104963 101354 105103
rect 123578 104963 123654 105103
rect 123878 104963 123954 105103
rect 146078 104963 146154 105103
rect 146578 104963 146654 105103
rect 168578 104963 168654 105103
rect 169478 104963 169554 105103
rect 190078 104963 190154 105103
rect 192178 104963 192254 105103
rect 208578 104963 208654 105103
rect 218678 104963 218754 105103
rect 11078 81828 11154 82103
rect 11193 81828 11269 82103
rect 33578 81828 33654 82103
rect 33696 81828 33772 82103
rect 56078 81828 56154 82103
rect 56203 81828 56279 82103
rect 78578 81828 78654 82103
rect 78728 81828 78804 82103
rect 101078 81828 101154 82103
rect 101278 81828 101354 82103
rect 123578 81828 123654 82103
rect 123878 81828 123954 82103
rect 146078 81828 146154 82103
rect 146578 81828 146654 82103
rect 168578 81828 168654 82103
rect 169478 81828 169554 82103
rect 190078 81828 190154 82103
rect 192178 81828 192254 82103
rect 208578 81828 208654 82103
rect 218678 81828 218754 82103
rect 11078 58628 11154 59103
rect 11193 58946 11269 59103
rect 11193 58633 11275 58946
rect 11193 58628 11269 58633
rect 33578 58628 33654 59103
rect 33696 58628 33772 59103
rect 56078 58628 56154 59103
rect 56203 58628 56279 59103
rect 78578 58628 78654 59103
rect 78728 58628 78804 59103
rect 101078 58628 101154 59103
rect 101278 58628 101354 59103
rect 123578 58628 123654 59103
rect 123878 58628 123954 59103
rect 146078 58628 146154 59103
rect 146578 58628 146654 59103
rect 168578 58628 168654 59103
rect 169478 58628 169554 59103
rect 190078 58628 190154 59103
rect 192178 58628 192254 59103
rect 208578 58628 208654 59103
rect 218678 58628 218754 59103
rect 11078 35428 11154 36103
rect 11193 35428 11269 36103
rect 33578 35428 33654 36103
rect 33696 35428 33772 36103
rect 56078 35428 56154 36103
rect 56203 35428 56279 36103
rect 78578 35428 78654 36103
rect 78728 35428 78804 36103
rect 101078 35428 101154 36103
rect 101278 35428 101354 36103
rect 123578 35428 123654 36103
rect 123878 35428 123954 36103
rect 146078 35428 146154 36103
rect 146578 35428 146654 36103
rect 168578 35428 168654 36103
rect 169478 35428 169554 36103
rect 190078 35428 190154 36103
rect 192178 35428 192254 36103
rect 208578 35428 208654 36103
rect 218678 35428 218754 36103
rect 11078 3128 11154 13103
rect 11193 3128 11269 13103
rect 33578 3128 33654 13103
rect 33696 3128 33772 13103
rect 56078 3128 56154 13103
rect 56203 3128 56279 13103
rect 78578 3128 78654 13103
rect 78728 3128 78804 13103
rect 101078 3128 101154 13103
rect 101278 3128 101354 13103
rect 123578 3128 123654 13103
rect 123878 3128 123954 13103
rect 146078 3128 146154 13103
rect 146578 3128 146654 13103
rect 168578 3128 168654 13103
rect 169478 3128 169554 13103
rect 190078 3128 190154 13103
rect 192178 3128 192254 13103
rect 208578 3128 208654 13103
rect 218678 3128 218754 13103
<< psubdiff >>
rect 10966 220103 11066 220116
rect 10966 220086 10979 220103
rect 11055 220086 11066 220103
rect 10966 220074 11066 220086
rect 33466 220103 33566 220116
rect 33466 220086 33479 220103
rect 33555 220086 33566 220103
rect 33466 220074 33566 220086
rect 55966 220103 56066 220116
rect 55966 220086 55979 220103
rect 56055 220086 56066 220103
rect 55966 220074 56066 220086
rect 78466 220103 78566 220116
rect 78466 220086 78479 220103
rect 78555 220086 78566 220103
rect 78466 220074 78566 220086
rect 100966 220103 101066 220116
rect 100966 220086 100979 220103
rect 101055 220086 101066 220103
rect 100966 220074 101066 220086
rect 123466 220103 123566 220116
rect 123466 220086 123479 220103
rect 123555 220086 123566 220103
rect 123466 220074 123566 220086
rect 145966 220103 146066 220116
rect 145966 220086 145979 220103
rect 146055 220086 146066 220103
rect 145966 220074 146066 220086
rect 168466 220103 168566 220116
rect 168466 220086 168479 220103
rect 168555 220086 168566 220103
rect 168466 220074 168566 220086
rect 189966 220103 190066 220116
rect 189966 220086 189979 220103
rect 190055 220086 190066 220103
rect 189966 220074 190066 220086
rect 192266 220074 192366 220116
rect 208466 220103 208566 220116
rect 208466 220086 208479 220103
rect 208555 220086 208566 220103
rect 208466 220074 208566 220086
rect 218766 220074 218866 220116
rect 10966 197103 11066 197116
rect 10966 197073 10979 197103
rect 11055 197073 11066 197103
rect 10966 197061 11066 197073
rect 33466 197103 33566 197116
rect 33466 197073 33479 197103
rect 33555 197073 33566 197103
rect 33466 197061 33566 197073
rect 55966 197103 56066 197116
rect 55966 197073 55979 197103
rect 56055 197073 56066 197103
rect 55966 197061 56066 197073
rect 78466 197103 78566 197116
rect 78466 197073 78479 197103
rect 78555 197073 78566 197103
rect 78466 197061 78566 197073
rect 100966 197103 101066 197116
rect 100966 197073 100979 197103
rect 101055 197073 101066 197103
rect 100966 197061 101066 197073
rect 123466 197103 123566 197116
rect 123466 197073 123479 197103
rect 123555 197073 123566 197103
rect 123466 197061 123566 197073
rect 145966 197103 146066 197116
rect 145966 197073 145979 197103
rect 146055 197073 146066 197103
rect 145966 197061 146066 197073
rect 168466 197103 168566 197116
rect 168466 197073 168479 197103
rect 168555 197073 168566 197103
rect 168466 197061 168566 197073
rect 189966 197103 190066 197116
rect 189966 197073 189979 197103
rect 190055 197073 190066 197103
rect 189966 197061 190066 197073
rect 192266 197061 192366 197116
rect 208466 197103 208566 197116
rect 208466 197073 208479 197103
rect 208555 197073 208566 197103
rect 208466 197061 208566 197073
rect 218766 197061 218866 197116
rect 10966 174103 11066 174116
rect 10966 174064 10979 174103
rect 11055 174064 11066 174103
rect 10966 174052 11066 174064
rect 33466 174103 33566 174116
rect 33466 174064 33479 174103
rect 33555 174064 33566 174103
rect 33466 174052 33566 174064
rect 55966 174103 56066 174116
rect 55966 174064 55979 174103
rect 56055 174064 56066 174103
rect 55966 174052 56066 174064
rect 78466 174103 78566 174116
rect 78466 174064 78479 174103
rect 78555 174064 78566 174103
rect 78466 174052 78566 174064
rect 100966 174103 101066 174116
rect 100966 174064 100979 174103
rect 101055 174064 101066 174103
rect 100966 174052 101066 174064
rect 123466 174103 123566 174116
rect 123466 174064 123479 174103
rect 123555 174064 123566 174103
rect 123466 174052 123566 174064
rect 145966 174103 146066 174116
rect 145966 174064 145979 174103
rect 146055 174064 146066 174103
rect 145966 174052 146066 174064
rect 168466 174103 168566 174116
rect 168466 174064 168479 174103
rect 168555 174064 168566 174103
rect 168466 174052 168566 174064
rect 189966 174103 190066 174116
rect 189966 174064 189979 174103
rect 190055 174064 190066 174103
rect 189966 174052 190066 174064
rect 192266 174052 192366 174116
rect 208466 174103 208566 174116
rect 208466 174064 208479 174103
rect 208555 174064 208566 174103
rect 208466 174052 208566 174064
rect 218766 174052 218866 174116
rect 10966 151103 11066 151116
rect 10966 151044 10979 151103
rect 11055 151044 11066 151103
rect 10966 151032 11066 151044
rect 33466 151103 33566 151116
rect 33466 151044 33479 151103
rect 33555 151044 33566 151103
rect 33466 151032 33566 151044
rect 55966 151103 56066 151116
rect 55966 151044 55979 151103
rect 56055 151044 56066 151103
rect 55966 151032 56066 151044
rect 78466 151103 78566 151116
rect 78466 151044 78479 151103
rect 78555 151044 78566 151103
rect 78466 151032 78566 151044
rect 100966 151103 101066 151116
rect 100966 151044 100979 151103
rect 101055 151044 101066 151103
rect 100966 151032 101066 151044
rect 123466 151103 123566 151116
rect 123466 151044 123479 151103
rect 123555 151044 123566 151103
rect 123466 151032 123566 151044
rect 145966 151103 146066 151116
rect 145966 151044 145979 151103
rect 146055 151044 146066 151103
rect 145966 151032 146066 151044
rect 168466 151103 168566 151116
rect 168466 151044 168479 151103
rect 168555 151044 168566 151103
rect 168466 151032 168566 151044
rect 189966 151103 190066 151116
rect 189966 151044 189979 151103
rect 190055 151044 190066 151103
rect 189966 151032 190066 151044
rect 192266 151032 192366 151116
rect 208466 151103 208566 151116
rect 208466 151044 208479 151103
rect 208555 151044 208566 151103
rect 208466 151032 208566 151044
rect 218766 151032 218866 151116
rect 10966 128103 11066 128116
rect 10966 128028 10979 128103
rect 11055 128028 11066 128103
rect 10966 128016 11066 128028
rect 33466 128103 33566 128116
rect 33466 128028 33479 128103
rect 33555 128028 33566 128103
rect 33466 128016 33566 128028
rect 55966 128103 56066 128116
rect 55966 128028 55979 128103
rect 56055 128028 56066 128103
rect 55966 128016 56066 128028
rect 78466 128103 78566 128116
rect 78466 128028 78479 128103
rect 78555 128028 78566 128103
rect 78466 128016 78566 128028
rect 100966 128103 101066 128116
rect 100966 128028 100979 128103
rect 101055 128028 101066 128103
rect 100966 128016 101066 128028
rect 123466 128103 123566 128116
rect 123466 128028 123479 128103
rect 123555 128028 123566 128103
rect 123466 128016 123566 128028
rect 145966 128103 146066 128116
rect 145966 128028 145979 128103
rect 146055 128028 146066 128103
rect 145966 128016 146066 128028
rect 168466 128103 168566 128116
rect 168466 128028 168479 128103
rect 168555 128028 168566 128103
rect 168466 128016 168566 128028
rect 189966 128103 190066 128116
rect 189966 128028 189979 128103
rect 190055 128028 190066 128103
rect 189966 128016 190066 128028
rect 192266 128016 192366 128116
rect 208466 128103 208566 128116
rect 208466 128028 208479 128103
rect 208555 128028 208566 128103
rect 208466 128016 208566 128028
rect 218766 128016 218866 128116
rect 10966 105103 11066 105116
rect 10966 104963 10979 105103
rect 11055 104963 11066 105103
rect 10966 104951 11066 104963
rect 33466 105103 33566 105116
rect 33466 104963 33479 105103
rect 33555 104963 33566 105103
rect 33466 104951 33566 104963
rect 55966 105103 56066 105116
rect 55966 104963 55979 105103
rect 56055 104963 56066 105103
rect 55966 104951 56066 104963
rect 78466 105103 78566 105116
rect 78466 104963 78479 105103
rect 78555 104963 78566 105103
rect 78466 104951 78566 104963
rect 100966 105103 101066 105116
rect 100966 104963 100979 105103
rect 101055 104963 101066 105103
rect 100966 104951 101066 104963
rect 123466 105103 123566 105116
rect 123466 104963 123479 105103
rect 123555 104963 123566 105103
rect 123466 104951 123566 104963
rect 145966 105103 146066 105116
rect 145966 104963 145979 105103
rect 146055 104963 146066 105103
rect 145966 104951 146066 104963
rect 168466 105103 168566 105116
rect 168466 104963 168479 105103
rect 168555 104963 168566 105103
rect 168466 104951 168566 104963
rect 189966 105103 190066 105116
rect 189966 104963 189979 105103
rect 190055 104963 190066 105103
rect 189966 104951 190066 104963
rect 192266 104951 192366 105116
rect 208466 105103 208566 105116
rect 208466 104963 208479 105103
rect 208555 104963 208566 105103
rect 208466 104951 208566 104963
rect 218766 104951 218866 105116
rect 10966 82103 11066 82116
rect 10966 81828 10979 82103
rect 11055 81828 11066 82103
rect 10966 81816 11066 81828
rect 33466 82103 33566 82116
rect 33466 81828 33479 82103
rect 33555 81828 33566 82103
rect 33466 81816 33566 81828
rect 55966 82103 56066 82116
rect 55966 81828 55979 82103
rect 56055 81828 56066 82103
rect 55966 81816 56066 81828
rect 78466 82103 78566 82116
rect 78466 81828 78479 82103
rect 78555 81828 78566 82103
rect 78466 81816 78566 81828
rect 100966 82103 101066 82116
rect 100966 81828 100979 82103
rect 101055 81828 101066 82103
rect 100966 81816 101066 81828
rect 123466 82103 123566 82116
rect 123466 81828 123479 82103
rect 123555 81828 123566 82103
rect 123466 81816 123566 81828
rect 145966 82103 146066 82116
rect 145966 81828 145979 82103
rect 146055 81828 146066 82103
rect 145966 81816 146066 81828
rect 168466 82103 168566 82116
rect 168466 81828 168479 82103
rect 168555 81828 168566 82103
rect 168466 81816 168566 81828
rect 189966 82103 190066 82116
rect 189966 81828 189979 82103
rect 190055 81828 190066 82103
rect 189966 81816 190066 81828
rect 192266 81816 192366 82116
rect 208466 82103 208566 82116
rect 208466 81828 208479 82103
rect 208555 81828 208566 82103
rect 208466 81816 208566 81828
rect 218766 81816 218866 82116
rect 10966 59103 11066 59116
rect 10966 58943 10979 59103
rect 10966 58633 10974 58943
rect 10966 58628 10979 58633
rect 11055 58628 11066 59103
rect 10966 58616 11066 58628
rect 33466 59103 33566 59116
rect 33466 58628 33479 59103
rect 33555 58628 33566 59103
rect 33466 58616 33566 58628
rect 55966 59103 56066 59116
rect 55966 58628 55979 59103
rect 56055 58628 56066 59103
rect 55966 58616 56066 58628
rect 78466 59103 78566 59116
rect 78466 58628 78479 59103
rect 78555 58628 78566 59103
rect 78466 58616 78566 58628
rect 100966 59103 101066 59116
rect 100966 58628 100979 59103
rect 101055 58628 101066 59103
rect 100966 58616 101066 58628
rect 123466 59103 123566 59116
rect 123466 58628 123479 59103
rect 123555 58628 123566 59103
rect 123466 58616 123566 58628
rect 145966 59103 146066 59116
rect 145966 58849 145979 59103
rect 145967 58628 145979 58849
rect 146055 58628 146066 59103
rect 145967 58616 146066 58628
rect 168466 59103 168566 59116
rect 168466 58628 168479 59103
rect 168555 58628 168566 59103
rect 168466 58616 168566 58628
rect 189966 59103 190066 59116
rect 189966 58628 189979 59103
rect 190055 58628 190066 59103
rect 189966 58616 190066 58628
rect 192266 58616 192366 59116
rect 208466 59103 208566 59116
rect 208466 58628 208479 59103
rect 208555 58628 208566 59103
rect 208466 58616 208566 58628
rect 218766 58616 218866 59116
rect 10966 36103 11066 36116
rect 10966 35428 10979 36103
rect 11055 35428 11066 36103
rect 10966 35416 11066 35428
rect 33466 36103 33566 36116
rect 33466 35428 33479 36103
rect 33555 35428 33566 36103
rect 33466 35416 33566 35428
rect 55966 36103 56066 36116
rect 55966 35428 55979 36103
rect 56055 35428 56066 36103
rect 55966 35416 56066 35428
rect 78466 36103 78566 36116
rect 78466 35428 78479 36103
rect 78555 35428 78566 36103
rect 78466 35416 78566 35428
rect 100966 36103 101066 36116
rect 100966 35428 100979 36103
rect 101055 35428 101066 36103
rect 100966 35416 101066 35428
rect 123466 36103 123566 36116
rect 123466 35428 123479 36103
rect 123555 35428 123566 36103
rect 123466 35416 123566 35428
rect 145966 36103 146066 36116
rect 145966 35428 145979 36103
rect 146055 35428 146066 36103
rect 145966 35416 146066 35428
rect 168466 36103 168566 36116
rect 168466 35428 168479 36103
rect 168555 35428 168566 36103
rect 168466 35416 168566 35428
rect 189966 36103 190066 36116
rect 189966 35428 189979 36103
rect 190055 35428 190066 36103
rect 189966 35416 190066 35428
rect 192266 35416 192366 36116
rect 208466 36103 208566 36116
rect 208466 35428 208479 36103
rect 208555 35428 208566 36103
rect 208466 35416 208566 35428
rect 218766 35416 218866 36116
rect 10966 13103 11066 13116
rect 10966 3128 10979 13103
rect 11055 3128 11066 13103
rect 10966 3116 11066 3128
rect 33466 13103 33566 13116
rect 33466 3128 33479 13103
rect 33555 3128 33566 13103
rect 33466 3116 33566 3128
rect 55966 13103 56066 13116
rect 55966 3128 55979 13103
rect 56055 3128 56066 13103
rect 55966 3116 56066 3128
rect 78466 13103 78566 13116
rect 78466 3128 78479 13103
rect 78555 3128 78566 13103
rect 78466 3116 78566 3128
rect 100966 13103 101066 13116
rect 100966 3128 100979 13103
rect 101055 3128 101066 13103
rect 100966 3116 101066 3128
rect 123466 13103 123566 13116
rect 123466 3128 123479 13103
rect 123555 3128 123566 13103
rect 123466 3116 123566 3128
rect 145966 13103 146066 13116
rect 145966 3128 145979 13103
rect 146055 3128 146066 13103
rect 145966 3116 146066 3128
rect 168466 13103 168566 13116
rect 168466 3128 168479 13103
rect 168555 3128 168566 13103
rect 168466 3116 168566 3128
rect 189966 13103 190066 13116
rect 189966 3128 189979 13103
rect 190055 3128 190066 13103
rect 189966 3116 190066 3128
rect 192266 3116 192366 13116
rect 208466 13103 208566 13116
rect 208466 3128 208479 13103
rect 208555 3128 208566 13103
rect 208466 3116 208566 3128
rect 218766 3116 218866 13116
<< psubdiffcont >>
rect 10979 220086 11055 220103
rect 33479 220086 33555 220103
rect 55979 220086 56055 220103
rect 78479 220086 78555 220103
rect 100979 220086 101055 220103
rect 123479 220086 123555 220103
rect 145979 220086 146055 220103
rect 168479 220086 168555 220103
rect 189979 220086 190055 220103
rect 208479 220086 208555 220103
rect 10979 197073 11055 197103
rect 33479 197073 33555 197103
rect 55979 197073 56055 197103
rect 78479 197073 78555 197103
rect 100979 197073 101055 197103
rect 123479 197073 123555 197103
rect 145979 197073 146055 197103
rect 168479 197073 168555 197103
rect 189979 197073 190055 197103
rect 208479 197073 208555 197103
rect 10979 174064 11055 174103
rect 33479 174064 33555 174103
rect 55979 174064 56055 174103
rect 78479 174064 78555 174103
rect 100979 174064 101055 174103
rect 123479 174064 123555 174103
rect 145979 174064 146055 174103
rect 168479 174064 168555 174103
rect 189979 174064 190055 174103
rect 208479 174064 208555 174103
rect 10979 151044 11055 151103
rect 33479 151044 33555 151103
rect 55979 151044 56055 151103
rect 78479 151044 78555 151103
rect 100979 151044 101055 151103
rect 123479 151044 123555 151103
rect 145979 151044 146055 151103
rect 168479 151044 168555 151103
rect 189979 151044 190055 151103
rect 208479 151044 208555 151103
rect 10979 128028 11055 128103
rect 33479 128028 33555 128103
rect 55979 128028 56055 128103
rect 78479 128028 78555 128103
rect 100979 128028 101055 128103
rect 123479 128028 123555 128103
rect 145979 128028 146055 128103
rect 168479 128028 168555 128103
rect 189979 128028 190055 128103
rect 208479 128028 208555 128103
rect 10979 104963 11055 105103
rect 33479 104963 33555 105103
rect 55979 104963 56055 105103
rect 78479 104963 78555 105103
rect 100979 104963 101055 105103
rect 123479 104963 123555 105103
rect 145979 104963 146055 105103
rect 168479 104963 168555 105103
rect 189979 104963 190055 105103
rect 208479 104963 208555 105103
rect 10979 81828 11055 82103
rect 33479 81828 33555 82103
rect 55979 81828 56055 82103
rect 78479 81828 78555 82103
rect 100979 81828 101055 82103
rect 123479 81828 123555 82103
rect 145979 81828 146055 82103
rect 168479 81828 168555 82103
rect 189979 81828 190055 82103
rect 208479 81828 208555 82103
rect 10979 58943 11055 59103
rect 10974 58633 11055 58943
rect 10979 58628 11055 58633
rect 33479 58628 33555 59103
rect 55979 58628 56055 59103
rect 78479 58628 78555 59103
rect 100979 58628 101055 59103
rect 123479 58628 123555 59103
rect 145979 58628 146055 59103
rect 168479 58628 168555 59103
rect 189979 58628 190055 59103
rect 208479 58628 208555 59103
rect 10979 35428 11055 36103
rect 33479 35428 33555 36103
rect 55979 35428 56055 36103
rect 78479 35428 78555 36103
rect 100979 35428 101055 36103
rect 123479 35428 123555 36103
rect 145979 35428 146055 36103
rect 168479 35428 168555 36103
rect 189979 35428 190055 36103
rect 208479 35428 208555 36103
rect 10979 3128 11055 13103
rect 33479 3128 33555 13103
rect 55979 3128 56055 13103
rect 78479 3128 78555 13103
rect 100979 3128 101055 13103
rect 123479 3128 123555 13103
rect 145979 3128 146055 13103
rect 168479 3128 168555 13103
rect 189979 3128 190055 13103
rect 208479 3128 208555 13103
<< poly >>
rect 11149 220183 11199 220191
rect 11149 220149 11157 220183
rect 11191 220149 11199 220183
rect 11149 220141 11199 220149
rect 33649 220183 33699 220191
rect 33649 220149 33657 220183
rect 33691 220149 33699 220183
rect 33649 220141 33699 220149
rect 56149 220183 56199 220191
rect 56149 220149 56157 220183
rect 56191 220149 56199 220183
rect 56149 220141 56199 220149
rect 78649 220183 78716 220191
rect 78649 220149 78657 220183
rect 78691 220149 78716 220183
rect 78649 220141 78716 220149
rect 101149 220183 101199 220191
rect 101149 220149 101157 220183
rect 101191 220149 101199 220183
rect 101149 220141 101199 220149
rect 123649 220183 123866 220191
rect 123649 220149 123657 220183
rect 123860 220149 123866 220183
rect 123649 220141 123866 220149
rect 146149 220183 146566 220191
rect 146149 220149 146157 220183
rect 146149 220148 146178 220149
rect 146552 220148 146566 220183
rect 146149 220141 146566 220148
rect 168649 220183 169462 220191
rect 168649 220149 168657 220183
rect 168649 220148 168680 220149
rect 169445 220148 169462 220183
rect 168649 220141 169462 220148
rect 190171 220184 192155 220191
rect 213649 220187 213699 220191
rect 190171 220150 190186 220184
rect 192127 220150 192155 220184
rect 190171 220149 191157 220150
rect 191191 220149 192155 220150
rect 190171 220141 192155 220149
rect 208669 220183 218659 220187
rect 208669 220178 213657 220183
rect 213691 220178 218659 220183
rect 208669 220148 208679 220178
rect 218645 220148 218659 220178
rect 11166 220116 11181 220141
rect 33666 220116 33685 220141
rect 56166 220116 56191 220141
rect 78666 220116 78716 220141
rect 101166 220116 101266 220141
rect 123666 220116 123866 220141
rect 146166 220116 146566 220141
rect 168666 220116 169466 220141
rect 190166 220116 192166 220141
rect 208669 220136 218659 220148
rect 208666 220134 218659 220136
rect 208666 220116 218666 220134
rect 11166 220059 11181 220074
rect 33666 220059 33685 220074
rect 56166 220059 56191 220074
rect 78666 220059 78716 220074
rect 101166 220059 101266 220074
rect 123666 220059 123866 220074
rect 146166 220059 146566 220074
rect 168666 220059 169466 220074
rect 190166 220059 192166 220074
rect 208666 220061 218666 220074
rect 213638 220059 218666 220061
rect 11149 197183 11199 197191
rect 11149 197149 11157 197183
rect 11191 197149 11199 197183
rect 11149 197141 11199 197149
rect 33649 197183 33699 197191
rect 33649 197149 33657 197183
rect 33691 197149 33699 197183
rect 33649 197141 33699 197149
rect 56149 197183 56199 197191
rect 56149 197149 56157 197183
rect 56191 197149 56199 197183
rect 56149 197141 56199 197149
rect 78649 197183 78716 197191
rect 78649 197149 78657 197183
rect 78691 197149 78716 197183
rect 78649 197141 78716 197149
rect 101149 197183 101199 197191
rect 101149 197149 101157 197183
rect 101191 197149 101199 197183
rect 101149 197141 101199 197149
rect 123649 197183 123866 197191
rect 123649 197149 123657 197183
rect 123860 197149 123866 197183
rect 123649 197141 123866 197149
rect 146149 197183 146566 197191
rect 146149 197149 146157 197183
rect 146149 197148 146178 197149
rect 146552 197148 146566 197183
rect 146149 197141 146566 197148
rect 168649 197183 169462 197191
rect 168649 197149 168657 197183
rect 168649 197148 168680 197149
rect 169445 197148 169462 197183
rect 168649 197141 169462 197148
rect 190171 197184 192155 197191
rect 213649 197187 213699 197191
rect 190171 197150 190186 197184
rect 192127 197150 192155 197184
rect 190171 197149 191157 197150
rect 191191 197149 192155 197150
rect 190171 197141 192155 197149
rect 208669 197183 218659 197187
rect 208669 197178 213657 197183
rect 213691 197178 218659 197183
rect 208669 197148 208679 197178
rect 218645 197148 218659 197178
rect 11166 197116 11181 197141
rect 33666 197116 33685 197141
rect 56166 197116 56191 197141
rect 78666 197116 78716 197141
rect 101166 197116 101266 197141
rect 123666 197116 123866 197141
rect 146166 197116 146566 197141
rect 168666 197116 169466 197141
rect 190166 197116 192166 197141
rect 208669 197136 218659 197148
rect 208666 197134 218659 197136
rect 208666 197116 218666 197134
rect 11166 197048 11181 197061
rect 33666 197048 33685 197061
rect 56166 197048 56191 197061
rect 78666 197048 78716 197061
rect 101166 197047 101266 197061
rect 123666 197047 123866 197061
rect 146166 197047 146566 197061
rect 168666 197048 169466 197061
rect 190166 197048 192166 197061
rect 208666 197048 218666 197061
rect 11149 174183 11199 174191
rect 11149 174149 11157 174183
rect 11191 174149 11199 174183
rect 11149 174141 11199 174149
rect 33649 174183 33699 174191
rect 33649 174149 33657 174183
rect 33691 174149 33699 174183
rect 33649 174141 33699 174149
rect 56149 174183 56199 174191
rect 56149 174149 56157 174183
rect 56191 174149 56199 174183
rect 56149 174141 56199 174149
rect 78649 174183 78716 174191
rect 78649 174149 78657 174183
rect 78691 174149 78716 174183
rect 78649 174141 78716 174149
rect 101149 174183 101199 174191
rect 101149 174149 101157 174183
rect 101191 174149 101199 174183
rect 101149 174141 101199 174149
rect 123649 174183 123866 174191
rect 123649 174149 123657 174183
rect 123860 174149 123866 174183
rect 123649 174141 123866 174149
rect 146149 174183 146566 174191
rect 146149 174149 146157 174183
rect 146149 174148 146178 174149
rect 146552 174148 146566 174183
rect 146149 174141 146566 174148
rect 168649 174183 169462 174191
rect 168649 174149 168657 174183
rect 168649 174148 168680 174149
rect 169445 174148 169462 174183
rect 168649 174141 169462 174148
rect 190171 174184 192155 174191
rect 213649 174187 213699 174191
rect 190171 174150 190186 174184
rect 192127 174150 192155 174184
rect 190171 174149 191157 174150
rect 191191 174149 192155 174150
rect 190171 174141 192155 174149
rect 208669 174183 218659 174187
rect 208669 174178 213657 174183
rect 213691 174178 218659 174183
rect 208669 174148 208679 174178
rect 218645 174148 218659 174178
rect 11166 174116 11181 174141
rect 33666 174116 33685 174141
rect 56166 174116 56191 174141
rect 78666 174116 78716 174141
rect 101166 174116 101266 174141
rect 123666 174116 123866 174141
rect 146166 174116 146566 174141
rect 168666 174116 169466 174141
rect 190166 174116 192166 174141
rect 208669 174136 218659 174148
rect 208666 174134 218659 174136
rect 208666 174116 218666 174134
rect 11166 174039 11181 174052
rect 33666 174036 33685 174052
rect 56166 174034 56191 174052
rect 78666 174032 78716 174052
rect 101166 174035 101266 174052
rect 123666 174036 123866 174052
rect 146166 174033 146566 174052
rect 168666 174039 169466 174052
rect 190166 174039 192166 174052
rect 208666 174039 218666 174052
rect 11149 151183 11199 151191
rect 11149 151149 11157 151183
rect 11191 151149 11199 151183
rect 11149 151141 11199 151149
rect 33649 151183 33699 151191
rect 33649 151149 33657 151183
rect 33691 151149 33699 151183
rect 33649 151141 33699 151149
rect 56149 151183 56199 151191
rect 56149 151149 56157 151183
rect 56191 151149 56199 151183
rect 56149 151141 56199 151149
rect 78649 151183 78716 151191
rect 78649 151149 78657 151183
rect 78691 151149 78716 151183
rect 78649 151141 78716 151149
rect 101149 151183 101199 151191
rect 101149 151149 101157 151183
rect 101191 151149 101199 151183
rect 101149 151141 101199 151149
rect 123649 151183 123866 151191
rect 123649 151149 123657 151183
rect 123860 151149 123866 151183
rect 123649 151141 123866 151149
rect 146149 151183 146566 151191
rect 146149 151149 146157 151183
rect 146149 151148 146178 151149
rect 146552 151148 146566 151183
rect 146149 151141 146566 151148
rect 168649 151183 169462 151191
rect 168649 151149 168657 151183
rect 168649 151148 168680 151149
rect 169445 151148 169462 151183
rect 168649 151141 169462 151148
rect 190171 151184 192155 151191
rect 213649 151187 213699 151191
rect 190171 151150 190186 151184
rect 192127 151150 192155 151184
rect 190171 151149 191157 151150
rect 191191 151149 192155 151150
rect 190171 151141 192155 151149
rect 208669 151183 218659 151187
rect 208669 151178 213657 151183
rect 213691 151178 218659 151183
rect 208669 151148 208679 151178
rect 218645 151148 218659 151178
rect 11166 151116 11181 151141
rect 33666 151116 33685 151141
rect 56166 151116 56191 151141
rect 78666 151116 78716 151141
rect 101166 151116 101266 151141
rect 123666 151116 123866 151141
rect 146166 151116 146566 151141
rect 168666 151116 169466 151141
rect 190166 151116 192166 151141
rect 208669 151136 218659 151148
rect 208666 151134 218659 151136
rect 208666 151116 218666 151134
rect 11166 151015 11181 151032
rect 33666 151008 33685 151032
rect 56166 151018 56191 151032
rect 78666 151015 78716 151032
rect 101166 151018 101266 151032
rect 123666 151006 123866 151032
rect 146166 151002 146566 151032
rect 168666 151012 169466 151032
rect 190166 151012 192166 151032
rect 208666 151017 218666 151032
rect 11149 128183 11199 128191
rect 11149 128149 11157 128183
rect 11191 128149 11199 128183
rect 11149 128141 11199 128149
rect 33649 128183 33699 128191
rect 33649 128149 33657 128183
rect 33691 128149 33699 128183
rect 33649 128141 33699 128149
rect 56149 128183 56199 128191
rect 56149 128149 56157 128183
rect 56191 128149 56199 128183
rect 56149 128141 56199 128149
rect 78649 128183 78716 128191
rect 78649 128149 78657 128183
rect 78691 128149 78716 128183
rect 78649 128141 78716 128149
rect 101149 128183 101199 128191
rect 101149 128149 101157 128183
rect 101191 128149 101199 128183
rect 101149 128141 101199 128149
rect 123649 128183 123866 128191
rect 123649 128149 123657 128183
rect 123860 128149 123866 128183
rect 123649 128141 123866 128149
rect 146149 128183 146566 128191
rect 146149 128149 146157 128183
rect 146149 128148 146178 128149
rect 146552 128148 146566 128183
rect 146149 128141 146566 128148
rect 168649 128183 169462 128191
rect 168649 128149 168657 128183
rect 168649 128148 168680 128149
rect 169445 128148 169462 128183
rect 168649 128141 169462 128148
rect 190171 128184 192155 128191
rect 213649 128187 213699 128191
rect 190171 128150 190186 128184
rect 192127 128150 192155 128184
rect 190171 128149 191157 128150
rect 191191 128149 192155 128150
rect 190171 128141 192155 128149
rect 208669 128183 218659 128187
rect 208669 128178 213657 128183
rect 213691 128178 218659 128183
rect 208669 128148 208679 128178
rect 218645 128148 218659 128178
rect 11166 128116 11181 128141
rect 33666 128116 33685 128141
rect 56166 128116 56191 128141
rect 78666 128116 78716 128141
rect 101166 128116 101266 128141
rect 123666 128116 123866 128141
rect 146166 128116 146566 128141
rect 168666 128116 169466 128141
rect 190166 128116 192166 128141
rect 208669 128136 218659 128148
rect 208666 128134 218659 128136
rect 208666 128116 218666 128134
rect 11166 128001 11181 128016
rect 33666 127997 33685 128016
rect 56166 128000 56191 128016
rect 78666 127991 78716 128016
rect 101166 127995 101266 128016
rect 123666 127995 123866 128016
rect 146166 127984 146566 128016
rect 168666 127987 169466 128016
rect 190166 127986 192166 128016
rect 208666 127990 218666 128016
rect 11149 105183 11199 105191
rect 11149 105149 11157 105183
rect 11191 105149 11199 105183
rect 11149 105141 11199 105149
rect 33649 105183 33699 105191
rect 33649 105149 33657 105183
rect 33691 105149 33699 105183
rect 33649 105141 33699 105149
rect 56149 105183 56199 105191
rect 56149 105149 56157 105183
rect 56191 105149 56199 105183
rect 56149 105141 56199 105149
rect 78649 105183 78716 105191
rect 78649 105149 78657 105183
rect 78691 105149 78716 105183
rect 78649 105141 78716 105149
rect 101149 105183 101199 105191
rect 101149 105149 101157 105183
rect 101191 105149 101199 105183
rect 101149 105141 101199 105149
rect 123649 105183 123866 105191
rect 123649 105149 123657 105183
rect 123860 105149 123866 105183
rect 123649 105141 123866 105149
rect 146149 105183 146566 105191
rect 146149 105149 146157 105183
rect 146149 105148 146178 105149
rect 146552 105148 146566 105183
rect 146149 105141 146566 105148
rect 168649 105183 169462 105191
rect 168649 105149 168657 105183
rect 168649 105148 168680 105149
rect 169445 105148 169462 105183
rect 168649 105141 169462 105148
rect 190171 105184 192155 105191
rect 213649 105187 213699 105191
rect 190171 105150 190186 105184
rect 192127 105150 192155 105184
rect 190171 105149 191157 105150
rect 191191 105149 192155 105150
rect 190171 105141 192155 105149
rect 208669 105183 218659 105187
rect 208669 105178 213657 105183
rect 213691 105178 218659 105183
rect 208669 105148 208679 105178
rect 218645 105148 218659 105178
rect 11166 105116 11181 105141
rect 33666 105116 33685 105141
rect 56166 105116 56191 105141
rect 78666 105116 78716 105141
rect 101166 105116 101266 105141
rect 123666 105116 123866 105141
rect 146166 105116 146566 105141
rect 168666 105116 169466 105141
rect 190166 105116 192166 105141
rect 208669 105136 218659 105148
rect 208666 105134 218659 105136
rect 208666 105116 218666 105134
rect 11166 104936 11181 104951
rect 33666 104936 33685 104951
rect 56166 104932 56191 104951
rect 78666 104931 78716 104951
rect 101166 104922 101266 104951
rect 123666 104917 123866 104951
rect 146166 104930 146566 104951
rect 168666 104929 169466 104951
rect 190166 104935 192166 104951
rect 208666 104936 218666 104951
rect 11149 82183 11199 82191
rect 11149 82149 11157 82183
rect 11191 82149 11199 82183
rect 11149 82141 11199 82149
rect 33649 82183 33699 82191
rect 33649 82149 33657 82183
rect 33691 82149 33699 82183
rect 33649 82141 33699 82149
rect 56149 82183 56199 82191
rect 56149 82149 56157 82183
rect 56191 82149 56199 82183
rect 56149 82141 56199 82149
rect 78649 82183 78716 82191
rect 78649 82149 78657 82183
rect 78691 82149 78716 82183
rect 78649 82141 78716 82149
rect 101149 82183 101199 82191
rect 101149 82149 101157 82183
rect 101191 82149 101199 82183
rect 101149 82141 101199 82149
rect 123649 82183 123866 82191
rect 123649 82149 123657 82183
rect 123860 82149 123866 82183
rect 123649 82141 123866 82149
rect 146149 82183 146566 82191
rect 146149 82149 146157 82183
rect 146149 82148 146178 82149
rect 146552 82148 146566 82183
rect 146149 82141 146566 82148
rect 168649 82183 169462 82191
rect 168649 82149 168657 82183
rect 168649 82148 168680 82149
rect 169445 82148 169462 82183
rect 168649 82141 169462 82148
rect 190171 82184 192155 82191
rect 213649 82187 213699 82191
rect 190171 82150 190186 82184
rect 192127 82150 192155 82184
rect 190171 82149 191157 82150
rect 191191 82149 192155 82150
rect 190171 82141 192155 82149
rect 208669 82183 218659 82187
rect 208669 82178 213657 82183
rect 213691 82178 218659 82183
rect 208669 82148 208679 82178
rect 218645 82148 218659 82178
rect 11166 82116 11181 82141
rect 33666 82116 33685 82141
rect 56166 82116 56191 82141
rect 78666 82116 78716 82141
rect 101166 82116 101266 82141
rect 123666 82116 123866 82141
rect 146166 82116 146566 82141
rect 168666 82116 169466 82141
rect 190166 82116 192166 82141
rect 208669 82136 218659 82148
rect 208666 82134 218659 82136
rect 208666 82116 218666 82134
rect 11166 81800 11181 81816
rect 33666 81798 33685 81816
rect 56166 81801 56191 81816
rect 78666 81798 78716 81816
rect 101166 81789 101266 81816
rect 123666 81798 123866 81816
rect 146166 81794 146566 81816
rect 168666 81797 169466 81816
rect 190166 81795 192166 81816
rect 208666 81795 218666 81816
rect 11149 59183 11199 59191
rect 11149 59149 11157 59183
rect 11191 59149 11199 59183
rect 11149 59141 11199 59149
rect 33649 59183 33699 59191
rect 33649 59149 33657 59183
rect 33691 59149 33699 59183
rect 33649 59141 33699 59149
rect 56149 59183 56199 59191
rect 56149 59149 56157 59183
rect 56191 59149 56199 59183
rect 56149 59141 56199 59149
rect 78649 59183 78716 59191
rect 78649 59149 78657 59183
rect 78691 59149 78716 59183
rect 78649 59141 78716 59149
rect 101149 59183 101199 59191
rect 101149 59149 101157 59183
rect 101191 59149 101199 59183
rect 101149 59141 101199 59149
rect 123649 59183 123866 59191
rect 123649 59149 123657 59183
rect 123860 59149 123866 59183
rect 123649 59141 123866 59149
rect 146149 59183 146566 59191
rect 146149 59149 146157 59183
rect 146149 59148 146178 59149
rect 146552 59148 146566 59183
rect 146149 59141 146566 59148
rect 168649 59183 169462 59191
rect 168649 59149 168657 59183
rect 168649 59148 168680 59149
rect 169445 59148 169462 59183
rect 168649 59141 169462 59148
rect 190171 59184 192155 59191
rect 213649 59187 213699 59191
rect 190171 59150 190186 59184
rect 192127 59150 192155 59184
rect 190171 59149 191157 59150
rect 191191 59149 192155 59150
rect 190171 59141 192155 59149
rect 208669 59183 218659 59187
rect 208669 59178 213657 59183
rect 213691 59178 218659 59183
rect 208669 59148 208679 59178
rect 218645 59148 218659 59178
rect 11166 59116 11181 59141
rect 33666 59116 33685 59141
rect 56166 59116 56191 59141
rect 78666 59116 78716 59141
rect 101166 59116 101266 59141
rect 123666 59116 123866 59141
rect 146166 59116 146566 59141
rect 168666 59116 169466 59141
rect 190166 59116 192166 59141
rect 208669 59136 218659 59148
rect 208666 59134 218659 59136
rect 208666 59116 218666 59134
rect 11166 58587 11181 58616
rect 33666 58588 33685 58616
rect 56166 58598 56191 58616
rect 78666 58594 78716 58616
rect 101166 58578 101266 58616
rect 123666 58578 123866 58616
rect 146166 58590 146566 58616
rect 168666 58598 169466 58616
rect 190166 58545 192166 58616
rect 208666 58597 218666 58616
rect 11149 36183 11199 36191
rect 11149 36149 11157 36183
rect 11191 36149 11199 36183
rect 11149 36141 11199 36149
rect 33649 36183 33699 36191
rect 33649 36149 33657 36183
rect 33691 36149 33699 36183
rect 33649 36141 33699 36149
rect 56149 36183 56199 36191
rect 56149 36149 56157 36183
rect 56191 36149 56199 36183
rect 56149 36141 56199 36149
rect 78649 36183 78716 36191
rect 78649 36149 78657 36183
rect 78691 36149 78716 36183
rect 78649 36141 78716 36149
rect 101149 36183 101199 36191
rect 101149 36149 101157 36183
rect 101191 36149 101199 36183
rect 101149 36141 101199 36149
rect 123649 36183 123866 36191
rect 123649 36149 123657 36183
rect 123860 36149 123866 36183
rect 123649 36141 123866 36149
rect 146149 36183 146566 36191
rect 146149 36149 146157 36183
rect 146149 36148 146178 36149
rect 146552 36148 146566 36183
rect 146149 36141 146566 36148
rect 168649 36183 169462 36191
rect 168649 36149 168657 36183
rect 168649 36148 168680 36149
rect 169445 36148 169462 36183
rect 168649 36141 169462 36148
rect 190171 36184 192155 36191
rect 213649 36187 213699 36191
rect 190171 36150 190186 36184
rect 192127 36150 192155 36184
rect 190171 36149 191157 36150
rect 191191 36149 192155 36150
rect 190171 36141 192155 36149
rect 208669 36183 218659 36187
rect 208669 36178 213657 36183
rect 213691 36178 218659 36183
rect 208669 36148 208679 36178
rect 218645 36148 218659 36178
rect 11166 36116 11181 36141
rect 33666 36116 33685 36141
rect 56166 36116 56191 36141
rect 78666 36116 78716 36141
rect 101166 36116 101266 36141
rect 123666 36116 123866 36141
rect 146166 36116 146566 36141
rect 168666 36116 169466 36141
rect 190166 36116 192166 36141
rect 208669 36136 218659 36148
rect 208666 36134 218659 36136
rect 208666 36116 218666 36134
rect 11166 35400 11181 35416
rect 33666 35397 33685 35416
rect 56166 35388 56191 35416
rect 78666 35386 78716 35416
rect 101166 35393 101266 35416
rect 123666 35391 123866 35416
rect 146166 35395 146566 35416
rect 168666 35388 169466 35416
rect 190166 35399 192166 35416
rect 208666 35382 218666 35416
rect 11149 13183 11199 13191
rect 11149 13149 11157 13183
rect 11191 13149 11199 13183
rect 11149 13141 11199 13149
rect 33649 13183 33699 13191
rect 33649 13149 33657 13183
rect 33691 13149 33699 13183
rect 33649 13141 33699 13149
rect 56149 13183 56199 13191
rect 56149 13149 56157 13183
rect 56191 13149 56199 13183
rect 56149 13141 56199 13149
rect 78649 13183 78716 13191
rect 78649 13149 78657 13183
rect 78691 13149 78716 13183
rect 78649 13141 78716 13149
rect 101149 13183 101199 13191
rect 101149 13149 101157 13183
rect 101191 13149 101199 13183
rect 101149 13141 101199 13149
rect 123649 13183 123866 13191
rect 123649 13149 123657 13183
rect 123860 13149 123866 13183
rect 123649 13141 123866 13149
rect 146149 13183 146566 13191
rect 146149 13149 146157 13183
rect 146149 13148 146178 13149
rect 146552 13148 146566 13183
rect 146149 13141 146566 13148
rect 168649 13183 169462 13191
rect 168649 13149 168657 13183
rect 168649 13148 168680 13149
rect 169445 13148 169462 13183
rect 168649 13141 169462 13148
rect 190171 13184 192155 13191
rect 213649 13187 213699 13191
rect 190171 13150 190186 13184
rect 192127 13150 192155 13184
rect 190171 13149 191157 13150
rect 191191 13149 192155 13150
rect 190171 13141 192155 13149
rect 208669 13183 218659 13187
rect 208669 13178 213657 13183
rect 213691 13178 218659 13183
rect 208669 13148 208679 13178
rect 218645 13148 218659 13178
rect 11166 13116 11181 13141
rect 33666 13116 33685 13141
rect 56166 13116 56191 13141
rect 78666 13116 78716 13141
rect 101166 13116 101266 13141
rect 123666 13116 123866 13141
rect 146166 13116 146566 13141
rect 168666 13116 169466 13141
rect 190166 13116 192166 13141
rect 208669 13136 218659 13148
rect 208666 13134 218659 13136
rect 208666 13116 218666 13134
rect 11166 3100 11181 3116
rect 33666 3097 33685 3116
rect 56166 3097 56191 3116
rect 78666 3084 78716 3116
rect 101166 3050 101266 3116
rect 123666 3058 123866 3116
rect 146166 3076 146566 3116
rect 168666 3091 169466 3116
rect 190166 3092 192166 3116
rect 208666 3090 218666 3116
<< polycont >>
rect 11157 220149 11191 220183
rect 33657 220149 33691 220183
rect 56157 220149 56191 220183
rect 78657 220149 78691 220183
rect 101157 220149 101191 220183
rect 123657 220149 123860 220183
rect 146157 220149 146552 220183
rect 146178 220148 146552 220149
rect 168657 220149 169445 220183
rect 168680 220148 169445 220149
rect 190186 220150 192127 220184
rect 191157 220149 191191 220150
rect 213657 220178 213691 220183
rect 208679 220148 218645 220178
rect 11157 197149 11191 197183
rect 33657 197149 33691 197183
rect 56157 197149 56191 197183
rect 78657 197149 78691 197183
rect 101157 197149 101191 197183
rect 123657 197149 123860 197183
rect 146157 197149 146552 197183
rect 146178 197148 146552 197149
rect 168657 197149 169445 197183
rect 168680 197148 169445 197149
rect 190186 197150 192127 197184
rect 191157 197149 191191 197150
rect 213657 197178 213691 197183
rect 208679 197148 218645 197178
rect 11157 174149 11191 174183
rect 33657 174149 33691 174183
rect 56157 174149 56191 174183
rect 78657 174149 78691 174183
rect 101157 174149 101191 174183
rect 123657 174149 123860 174183
rect 146157 174149 146552 174183
rect 146178 174148 146552 174149
rect 168657 174149 169445 174183
rect 168680 174148 169445 174149
rect 190186 174150 192127 174184
rect 191157 174149 191191 174150
rect 213657 174178 213691 174183
rect 208679 174148 218645 174178
rect 11157 151149 11191 151183
rect 33657 151149 33691 151183
rect 56157 151149 56191 151183
rect 78657 151149 78691 151183
rect 101157 151149 101191 151183
rect 123657 151149 123860 151183
rect 146157 151149 146552 151183
rect 146178 151148 146552 151149
rect 168657 151149 169445 151183
rect 168680 151148 169445 151149
rect 190186 151150 192127 151184
rect 191157 151149 191191 151150
rect 213657 151178 213691 151183
rect 208679 151148 218645 151178
rect 11157 128149 11191 128183
rect 33657 128149 33691 128183
rect 56157 128149 56191 128183
rect 78657 128149 78691 128183
rect 101157 128149 101191 128183
rect 123657 128149 123860 128183
rect 146157 128149 146552 128183
rect 146178 128148 146552 128149
rect 168657 128149 169445 128183
rect 168680 128148 169445 128149
rect 190186 128150 192127 128184
rect 191157 128149 191191 128150
rect 213657 128178 213691 128183
rect 208679 128148 218645 128178
rect 11157 105149 11191 105183
rect 33657 105149 33691 105183
rect 56157 105149 56191 105183
rect 78657 105149 78691 105183
rect 101157 105149 101191 105183
rect 123657 105149 123860 105183
rect 146157 105149 146552 105183
rect 146178 105148 146552 105149
rect 168657 105149 169445 105183
rect 168680 105148 169445 105149
rect 190186 105150 192127 105184
rect 191157 105149 191191 105150
rect 213657 105178 213691 105183
rect 208679 105148 218645 105178
rect 11157 82149 11191 82183
rect 33657 82149 33691 82183
rect 56157 82149 56191 82183
rect 78657 82149 78691 82183
rect 101157 82149 101191 82183
rect 123657 82149 123860 82183
rect 146157 82149 146552 82183
rect 146178 82148 146552 82149
rect 168657 82149 169445 82183
rect 168680 82148 169445 82149
rect 190186 82150 192127 82184
rect 191157 82149 191191 82150
rect 213657 82178 213691 82183
rect 208679 82148 218645 82178
rect 11157 59149 11191 59183
rect 33657 59149 33691 59183
rect 56157 59149 56191 59183
rect 78657 59149 78691 59183
rect 101157 59149 101191 59183
rect 123657 59149 123860 59183
rect 146157 59149 146552 59183
rect 146178 59148 146552 59149
rect 168657 59149 169445 59183
rect 168680 59148 169445 59149
rect 190186 59150 192127 59184
rect 191157 59149 191191 59150
rect 213657 59178 213691 59183
rect 208679 59148 218645 59178
rect 11157 36149 11191 36183
rect 33657 36149 33691 36183
rect 56157 36149 56191 36183
rect 78657 36149 78691 36183
rect 101157 36149 101191 36183
rect 123657 36149 123860 36183
rect 146157 36149 146552 36183
rect 146178 36148 146552 36149
rect 168657 36149 169445 36183
rect 168680 36148 169445 36149
rect 190186 36150 192127 36184
rect 191157 36149 191191 36150
rect 213657 36178 213691 36183
rect 208679 36148 218645 36178
rect 11157 13149 11191 13183
rect 33657 13149 33691 13183
rect 56157 13149 56191 13183
rect 78657 13149 78691 13183
rect 101157 13149 101191 13183
rect 123657 13149 123860 13183
rect 146157 13149 146552 13183
rect 146178 13148 146552 13149
rect 168657 13149 169445 13183
rect 168680 13148 169445 13149
rect 190186 13150 192127 13184
rect 191157 13149 191191 13150
rect 213657 13178 213691 13183
rect 208679 13148 218645 13178
<< locali >>
rect 11149 220183 11199 220191
rect 11149 220149 11157 220183
rect 11191 220149 11199 220183
rect 11149 220141 11199 220149
rect 33649 220183 33699 220191
rect 33649 220149 33657 220183
rect 33691 220149 33699 220183
rect 33649 220141 33699 220149
rect 56149 220183 56199 220191
rect 56149 220149 56157 220183
rect 56191 220149 56199 220183
rect 56149 220141 56199 220149
rect 78649 220183 78716 220191
rect 78649 220149 78657 220183
rect 78691 220149 78716 220183
rect 78649 220141 78716 220149
rect 101149 220183 101199 220191
rect 101149 220149 101157 220183
rect 101191 220149 101199 220183
rect 101149 220141 101199 220149
rect 123649 220183 123866 220191
rect 123649 220149 123657 220183
rect 123860 220149 123866 220183
rect 123649 220141 123866 220149
rect 146149 220183 146566 220191
rect 146149 220149 146157 220183
rect 146149 220148 146178 220149
rect 146552 220148 146566 220183
rect 146149 220141 146566 220148
rect 168649 220183 169463 220191
rect 168649 220149 168657 220183
rect 168649 220148 168680 220149
rect 169445 220148 169463 220183
rect 168649 220141 169463 220148
rect 190176 220184 192154 220191
rect 213649 220186 213699 220191
rect 190176 220150 190186 220184
rect 192127 220150 192154 220184
rect 190176 220149 191157 220150
rect 191191 220149 192154 220150
rect 190176 220146 192154 220149
rect 208670 220183 218658 220186
rect 208670 220178 213657 220183
rect 213691 220178 218658 220183
rect 208670 220148 208679 220178
rect 218645 220148 218658 220178
rect 191149 220141 191199 220146
rect 208670 220140 218658 220148
rect 10968 220103 11056 220114
rect 10968 220086 10974 220103
rect 11055 220086 11056 220103
rect 10968 220076 11056 220086
rect 11076 220103 11164 220114
rect 11076 220086 11078 220103
rect 11154 220086 11164 220103
rect 11076 220076 11164 220086
rect 11183 220103 11279 220114
rect 11183 220086 11193 220103
rect 11274 220086 11279 220103
rect 11183 220076 11279 220086
rect 33468 220103 33556 220114
rect 33468 220086 33474 220103
rect 33555 220086 33556 220103
rect 33468 220076 33556 220086
rect 33576 220103 33664 220114
rect 33576 220086 33578 220103
rect 33654 220086 33664 220103
rect 33576 220076 33664 220086
rect 33686 220103 33782 220114
rect 33686 220086 33696 220103
rect 33777 220086 33782 220103
rect 33686 220076 33782 220086
rect 55968 220103 56056 220114
rect 55968 220086 55974 220103
rect 56055 220086 56056 220103
rect 55968 220076 56056 220086
rect 56076 220103 56164 220114
rect 56076 220086 56078 220103
rect 56154 220086 56164 220103
rect 56076 220076 56164 220086
rect 56193 220103 56289 220114
rect 56193 220086 56203 220103
rect 56284 220086 56289 220103
rect 56193 220076 56289 220086
rect 78468 220103 78556 220114
rect 78468 220086 78474 220103
rect 78555 220086 78556 220103
rect 78468 220076 78556 220086
rect 78576 220103 78664 220114
rect 78576 220086 78578 220103
rect 78654 220086 78664 220103
rect 78576 220076 78664 220086
rect 78718 220103 78814 220114
rect 78718 220086 78728 220103
rect 78809 220086 78814 220103
rect 78718 220076 78814 220086
rect 100968 220103 101056 220114
rect 100968 220086 100974 220103
rect 101055 220086 101056 220103
rect 100968 220076 101056 220086
rect 101076 220103 101164 220114
rect 101076 220086 101078 220103
rect 101154 220086 101164 220103
rect 101076 220076 101164 220086
rect 101268 220103 101364 220114
rect 101268 220086 101278 220103
rect 101359 220086 101364 220103
rect 101268 220076 101364 220086
rect 123468 220103 123556 220114
rect 123468 220086 123474 220103
rect 123555 220086 123556 220103
rect 123468 220076 123556 220086
rect 123576 220103 123664 220114
rect 123576 220086 123578 220103
rect 123654 220086 123664 220103
rect 123576 220076 123664 220086
rect 123868 220103 123964 220114
rect 123868 220086 123878 220103
rect 123959 220086 123964 220103
rect 123868 220076 123964 220086
rect 145968 220103 146056 220114
rect 145968 220086 145974 220103
rect 146055 220086 146056 220103
rect 145968 220076 146056 220086
rect 146076 220103 146164 220114
rect 146076 220086 146078 220103
rect 146154 220086 146164 220103
rect 146076 220076 146164 220086
rect 146568 220103 146664 220114
rect 146568 220086 146578 220103
rect 146659 220086 146664 220103
rect 146568 220076 146664 220086
rect 168468 220103 168556 220114
rect 168468 220086 168474 220103
rect 168555 220086 168556 220103
rect 168468 220076 168556 220086
rect 168576 220103 168664 220114
rect 168576 220086 168578 220103
rect 168654 220086 168664 220103
rect 168576 220076 168664 220086
rect 169468 220103 169564 220114
rect 169468 220086 169478 220103
rect 169559 220086 169564 220103
rect 169468 220076 169564 220086
rect 189968 220103 190056 220114
rect 189968 220086 189974 220103
rect 190055 220086 190056 220103
rect 189968 220076 190056 220086
rect 190076 220103 190164 220114
rect 190076 220086 190078 220103
rect 190154 220086 190164 220103
rect 190076 220076 190164 220086
rect 192168 220103 192265 220114
rect 192168 220086 192178 220103
rect 192259 220086 192265 220103
rect 192168 220076 192265 220086
rect 208468 220103 208556 220114
rect 208468 220086 208474 220103
rect 208555 220086 208556 220103
rect 208468 220076 208556 220086
rect 208576 220103 208664 220114
rect 208576 220086 208578 220103
rect 208654 220086 208664 220103
rect 208576 220076 208664 220086
rect 218668 220103 218775 220114
rect 218668 220086 218678 220103
rect 218759 220086 218775 220103
rect 218668 220076 218775 220086
rect 11149 197183 11199 197191
rect 11149 197149 11157 197183
rect 11191 197149 11199 197183
rect 11149 197141 11199 197149
rect 33649 197183 33699 197191
rect 33649 197149 33657 197183
rect 33691 197149 33699 197183
rect 33649 197141 33699 197149
rect 56149 197183 56199 197191
rect 56149 197149 56157 197183
rect 56191 197149 56199 197183
rect 56149 197141 56199 197149
rect 78649 197183 78716 197191
rect 78649 197149 78657 197183
rect 78691 197149 78716 197183
rect 78649 197141 78716 197149
rect 101149 197183 101199 197191
rect 101149 197149 101157 197183
rect 101191 197149 101199 197183
rect 101149 197141 101199 197149
rect 123649 197183 123866 197191
rect 123649 197149 123657 197183
rect 123860 197149 123866 197183
rect 123649 197141 123866 197149
rect 146149 197183 146566 197191
rect 146149 197149 146157 197183
rect 146149 197148 146178 197149
rect 146552 197148 146566 197183
rect 146149 197141 146566 197148
rect 168649 197183 169463 197191
rect 168649 197149 168657 197183
rect 168649 197148 168680 197149
rect 169445 197148 169463 197183
rect 168649 197141 169463 197148
rect 190176 197184 192154 197191
rect 213649 197186 213699 197191
rect 190176 197150 190186 197184
rect 192127 197150 192154 197184
rect 190176 197149 191157 197150
rect 191191 197149 192154 197150
rect 190176 197146 192154 197149
rect 208670 197183 218658 197186
rect 208670 197178 213657 197183
rect 213691 197178 218658 197183
rect 208670 197148 208679 197178
rect 218645 197148 218658 197178
rect 191149 197141 191199 197146
rect 208670 197140 218658 197148
rect 10968 197103 11056 197114
rect 10968 197073 10974 197103
rect 11055 197073 11056 197103
rect 10968 197063 11056 197073
rect 11076 197103 11164 197114
rect 11076 197073 11078 197103
rect 11154 197073 11164 197103
rect 11076 197063 11164 197073
rect 11183 197103 11279 197114
rect 11183 197073 11193 197103
rect 11274 197073 11279 197103
rect 11183 197063 11279 197073
rect 33468 197103 33556 197114
rect 33468 197073 33474 197103
rect 33555 197073 33556 197103
rect 33468 197063 33556 197073
rect 33576 197103 33664 197114
rect 33576 197073 33578 197103
rect 33654 197073 33664 197103
rect 33576 197063 33664 197073
rect 33686 197103 33782 197114
rect 33686 197073 33696 197103
rect 33777 197073 33782 197103
rect 33686 197063 33782 197073
rect 55968 197103 56056 197114
rect 55968 197073 55974 197103
rect 56055 197073 56056 197103
rect 55968 197063 56056 197073
rect 56076 197103 56164 197114
rect 56076 197073 56078 197103
rect 56154 197073 56164 197103
rect 56076 197063 56164 197073
rect 56193 197103 56289 197114
rect 56193 197073 56203 197103
rect 56284 197073 56289 197103
rect 56193 197063 56289 197073
rect 78468 197103 78556 197114
rect 78468 197073 78474 197103
rect 78555 197073 78556 197103
rect 78468 197063 78556 197073
rect 78576 197103 78664 197114
rect 78576 197073 78578 197103
rect 78654 197073 78664 197103
rect 78576 197063 78664 197073
rect 78718 197103 78814 197114
rect 78718 197073 78728 197103
rect 78809 197073 78814 197103
rect 78718 197063 78814 197073
rect 100968 197103 101056 197114
rect 100968 197073 100974 197103
rect 101055 197073 101056 197103
rect 100968 197063 101056 197073
rect 101076 197103 101164 197114
rect 101076 197073 101078 197103
rect 101154 197073 101164 197103
rect 101076 197063 101164 197073
rect 101268 197103 101364 197114
rect 101268 197073 101278 197103
rect 101359 197073 101364 197103
rect 101268 197063 101364 197073
rect 123468 197103 123556 197114
rect 123468 197073 123474 197103
rect 123555 197073 123556 197103
rect 123468 197063 123556 197073
rect 123576 197103 123664 197114
rect 123576 197073 123578 197103
rect 123654 197073 123664 197103
rect 123576 197063 123664 197073
rect 123868 197103 123964 197114
rect 123868 197073 123878 197103
rect 123959 197073 123964 197103
rect 123868 197063 123964 197073
rect 145968 197103 146056 197114
rect 145968 197073 145974 197103
rect 146055 197073 146056 197103
rect 145968 197063 146056 197073
rect 146076 197103 146164 197114
rect 146076 197073 146078 197103
rect 146154 197073 146164 197103
rect 146076 197063 146164 197073
rect 146568 197103 146664 197114
rect 146568 197073 146578 197103
rect 146659 197073 146664 197103
rect 146568 197063 146664 197073
rect 168468 197103 168556 197114
rect 168468 197073 168474 197103
rect 168555 197073 168556 197103
rect 168468 197063 168556 197073
rect 168576 197103 168664 197114
rect 168576 197073 168578 197103
rect 168654 197073 168664 197103
rect 168576 197063 168664 197073
rect 169468 197103 169564 197114
rect 169468 197073 169478 197103
rect 169559 197073 169564 197103
rect 169468 197063 169564 197073
rect 189968 197103 190056 197114
rect 189968 197073 189974 197103
rect 190055 197073 190056 197103
rect 189968 197063 190056 197073
rect 190076 197103 190164 197114
rect 190076 197073 190078 197103
rect 190154 197073 190164 197103
rect 190076 197063 190164 197073
rect 192168 197103 192270 197114
rect 192168 197073 192178 197103
rect 192259 197073 192270 197103
rect 192168 197063 192270 197073
rect 208468 197103 208556 197114
rect 208468 197073 208474 197103
rect 208555 197073 208556 197103
rect 208468 197063 208556 197073
rect 208576 197103 208664 197114
rect 208576 197073 208578 197103
rect 208654 197073 208664 197103
rect 208576 197063 208664 197073
rect 218668 197103 218770 197114
rect 218668 197073 218678 197103
rect 218759 197073 218770 197103
rect 218668 197063 218770 197073
rect 11149 174183 11199 174191
rect 11149 174149 11157 174183
rect 11191 174149 11199 174183
rect 11149 174141 11199 174149
rect 33649 174183 33699 174191
rect 33649 174149 33657 174183
rect 33691 174149 33699 174183
rect 33649 174141 33699 174149
rect 56149 174183 56199 174191
rect 56149 174149 56157 174183
rect 56191 174149 56199 174183
rect 56149 174141 56199 174149
rect 78649 174183 78716 174191
rect 78649 174149 78657 174183
rect 78691 174149 78716 174183
rect 78649 174141 78716 174149
rect 101149 174183 101199 174191
rect 101149 174149 101157 174183
rect 101191 174149 101199 174183
rect 101149 174141 101199 174149
rect 123649 174183 123866 174191
rect 123649 174149 123657 174183
rect 123860 174149 123866 174183
rect 123649 174141 123866 174149
rect 146149 174183 146566 174191
rect 146149 174149 146157 174183
rect 146149 174148 146178 174149
rect 146552 174148 146566 174183
rect 146149 174141 146566 174148
rect 168649 174183 169463 174191
rect 168649 174149 168657 174183
rect 168649 174148 168680 174149
rect 169445 174148 169463 174183
rect 168649 174141 169463 174148
rect 190176 174184 192154 174191
rect 213649 174186 213699 174191
rect 190176 174150 190186 174184
rect 192127 174150 192154 174184
rect 190176 174149 191157 174150
rect 191191 174149 192154 174150
rect 190176 174146 192154 174149
rect 208670 174183 218658 174186
rect 208670 174178 213657 174183
rect 213691 174178 218658 174183
rect 208670 174148 208679 174178
rect 218645 174148 218658 174178
rect 191149 174141 191199 174146
rect 208670 174140 218658 174148
rect 10968 174103 11056 174114
rect 10968 174064 10974 174103
rect 11055 174064 11056 174103
rect 10968 174054 11056 174064
rect 11076 174103 11164 174114
rect 11076 174064 11078 174103
rect 11154 174064 11164 174103
rect 11076 174054 11164 174064
rect 11183 174103 11279 174114
rect 11183 174064 11193 174103
rect 11274 174064 11279 174103
rect 11183 174054 11279 174064
rect 33468 174103 33556 174114
rect 33468 174064 33474 174103
rect 33555 174064 33556 174103
rect 33468 174054 33556 174064
rect 33576 174103 33664 174114
rect 33576 174064 33578 174103
rect 33654 174064 33664 174103
rect 33576 174054 33664 174064
rect 33686 174103 33782 174114
rect 33686 174064 33696 174103
rect 33777 174064 33782 174103
rect 33686 174054 33782 174064
rect 55968 174103 56056 174114
rect 55968 174064 55974 174103
rect 56055 174064 56056 174103
rect 55968 174054 56056 174064
rect 56076 174103 56164 174114
rect 56076 174064 56078 174103
rect 56154 174064 56164 174103
rect 56076 174054 56164 174064
rect 56193 174103 56289 174114
rect 56193 174064 56203 174103
rect 56284 174064 56289 174103
rect 56193 174054 56289 174064
rect 78468 174103 78556 174114
rect 78468 174064 78474 174103
rect 78555 174064 78556 174103
rect 78468 174054 78556 174064
rect 78576 174103 78664 174114
rect 78576 174064 78578 174103
rect 78654 174064 78664 174103
rect 78576 174054 78664 174064
rect 78718 174103 78814 174114
rect 78718 174064 78728 174103
rect 78809 174064 78814 174103
rect 78718 174054 78814 174064
rect 100968 174103 101056 174114
rect 100968 174064 100974 174103
rect 101055 174064 101056 174103
rect 100968 174054 101056 174064
rect 101076 174103 101164 174114
rect 101076 174064 101078 174103
rect 101154 174064 101164 174103
rect 101076 174054 101164 174064
rect 101268 174103 101364 174114
rect 101268 174064 101278 174103
rect 101359 174064 101364 174103
rect 101268 174054 101364 174064
rect 123468 174103 123556 174114
rect 123468 174064 123474 174103
rect 123555 174064 123556 174103
rect 123468 174054 123556 174064
rect 123576 174103 123664 174114
rect 123576 174064 123578 174103
rect 123654 174064 123664 174103
rect 123576 174054 123664 174064
rect 123868 174103 123964 174114
rect 123868 174064 123878 174103
rect 123959 174064 123964 174103
rect 123868 174054 123964 174064
rect 145968 174103 146056 174114
rect 145968 174064 145974 174103
rect 146055 174064 146056 174103
rect 145968 174054 146056 174064
rect 146076 174103 146164 174114
rect 146076 174064 146078 174103
rect 146154 174064 146164 174103
rect 146076 174054 146164 174064
rect 146568 174103 146664 174114
rect 146568 174064 146578 174103
rect 146659 174064 146664 174103
rect 146568 174054 146664 174064
rect 168468 174103 168556 174114
rect 168468 174064 168474 174103
rect 168555 174064 168556 174103
rect 168468 174054 168556 174064
rect 168576 174103 168664 174114
rect 168576 174064 168578 174103
rect 168654 174064 168664 174103
rect 168576 174054 168664 174064
rect 169468 174103 169564 174114
rect 169468 174064 169478 174103
rect 169559 174064 169564 174103
rect 169468 174054 169564 174064
rect 189968 174103 190056 174114
rect 189968 174064 189974 174103
rect 190055 174064 190056 174103
rect 189968 174054 190056 174064
rect 190076 174103 190164 174114
rect 190076 174064 190078 174103
rect 190154 174064 190164 174103
rect 190076 174054 190164 174064
rect 192168 174103 192265 174114
rect 192168 174064 192178 174103
rect 192259 174064 192265 174103
rect 192168 174054 192265 174064
rect 208468 174103 208556 174114
rect 208468 174064 208474 174103
rect 208555 174064 208556 174103
rect 208468 174054 208556 174064
rect 208576 174103 208664 174114
rect 208576 174064 208578 174103
rect 208654 174064 208664 174103
rect 208576 174054 208664 174064
rect 218668 174103 218770 174114
rect 218668 174064 218678 174103
rect 218759 174064 218770 174103
rect 218668 174054 218770 174064
rect 11149 151183 11199 151191
rect 11149 151149 11157 151183
rect 11191 151149 11199 151183
rect 11149 151141 11199 151149
rect 33649 151183 33699 151191
rect 33649 151149 33657 151183
rect 33691 151149 33699 151183
rect 33649 151141 33699 151149
rect 56149 151183 56199 151191
rect 56149 151149 56157 151183
rect 56191 151149 56199 151183
rect 56149 151141 56199 151149
rect 78649 151183 78716 151191
rect 78649 151149 78657 151183
rect 78691 151149 78716 151183
rect 78649 151141 78716 151149
rect 101149 151183 101199 151191
rect 101149 151149 101157 151183
rect 101191 151149 101199 151183
rect 101149 151141 101199 151149
rect 123649 151183 123866 151191
rect 123649 151149 123657 151183
rect 123860 151149 123866 151183
rect 123649 151141 123866 151149
rect 146149 151183 146566 151191
rect 146149 151149 146157 151183
rect 146149 151148 146178 151149
rect 146552 151148 146566 151183
rect 146149 151141 146566 151148
rect 168649 151183 169463 151191
rect 168649 151149 168657 151183
rect 168649 151148 168680 151149
rect 169445 151148 169463 151183
rect 168649 151141 169463 151148
rect 190176 151184 192154 151191
rect 213649 151186 213699 151191
rect 190176 151150 190186 151184
rect 192127 151150 192154 151184
rect 190176 151149 191157 151150
rect 191191 151149 192154 151150
rect 190176 151146 192154 151149
rect 208670 151183 218658 151186
rect 208670 151178 213657 151183
rect 213691 151178 218658 151183
rect 208670 151148 208679 151178
rect 218645 151148 218658 151178
rect 191149 151141 191199 151146
rect 208670 151140 218658 151148
rect 10968 151103 11056 151114
rect 10968 151044 10974 151103
rect 11055 151044 11056 151103
rect 10968 151034 11056 151044
rect 11076 151103 11164 151114
rect 11076 151044 11078 151103
rect 11154 151044 11164 151103
rect 11076 151034 11164 151044
rect 11183 151103 11279 151114
rect 11183 151044 11193 151103
rect 11274 151044 11279 151103
rect 11183 151034 11279 151044
rect 33468 151103 33556 151114
rect 33468 151044 33474 151103
rect 33555 151044 33556 151103
rect 33468 151034 33556 151044
rect 33576 151103 33664 151114
rect 33576 151044 33578 151103
rect 33654 151044 33664 151103
rect 33576 151034 33664 151044
rect 33686 151103 33782 151114
rect 33686 151044 33696 151103
rect 33777 151044 33782 151103
rect 33686 151034 33782 151044
rect 55968 151103 56056 151114
rect 55968 151044 55974 151103
rect 56055 151044 56056 151103
rect 55968 151034 56056 151044
rect 56076 151103 56164 151114
rect 56076 151044 56078 151103
rect 56154 151044 56164 151103
rect 56076 151034 56164 151044
rect 56193 151103 56289 151114
rect 56193 151044 56203 151103
rect 56284 151044 56289 151103
rect 56193 151034 56289 151044
rect 78468 151103 78556 151114
rect 78468 151044 78474 151103
rect 78555 151044 78556 151103
rect 78468 151034 78556 151044
rect 78576 151103 78664 151114
rect 78576 151044 78578 151103
rect 78654 151044 78664 151103
rect 78576 151034 78664 151044
rect 78718 151103 78814 151114
rect 78718 151044 78728 151103
rect 78809 151044 78814 151103
rect 78718 151034 78814 151044
rect 100968 151103 101056 151114
rect 100968 151044 100974 151103
rect 101055 151044 101056 151103
rect 100968 151034 101056 151044
rect 101076 151103 101164 151114
rect 101076 151044 101078 151103
rect 101154 151044 101164 151103
rect 101076 151034 101164 151044
rect 101268 151103 101364 151114
rect 101268 151044 101278 151103
rect 101359 151044 101364 151103
rect 101268 151034 101364 151044
rect 123468 151103 123556 151114
rect 123468 151044 123474 151103
rect 123555 151044 123556 151103
rect 123468 151034 123556 151044
rect 123576 151103 123664 151114
rect 123576 151044 123578 151103
rect 123654 151044 123664 151103
rect 123576 151034 123664 151044
rect 123868 151103 123964 151114
rect 123868 151044 123878 151103
rect 123959 151044 123964 151103
rect 123868 151034 123964 151044
rect 145968 151103 146056 151114
rect 145968 151044 145974 151103
rect 146055 151044 146056 151103
rect 145968 151034 146056 151044
rect 146076 151103 146164 151114
rect 146076 151044 146078 151103
rect 146154 151044 146164 151103
rect 146076 151034 146164 151044
rect 146568 151103 146664 151114
rect 146568 151044 146578 151103
rect 146659 151044 146664 151103
rect 146568 151034 146664 151044
rect 168468 151103 168556 151114
rect 168468 151044 168474 151103
rect 168555 151044 168556 151103
rect 168468 151034 168556 151044
rect 168576 151103 168664 151114
rect 168576 151044 168578 151103
rect 168654 151044 168664 151103
rect 168576 151034 168664 151044
rect 169468 151103 169564 151114
rect 169468 151044 169478 151103
rect 169559 151044 169564 151103
rect 169468 151034 169564 151044
rect 189968 151103 190056 151114
rect 189968 151044 189974 151103
rect 190055 151044 190056 151103
rect 189968 151034 190056 151044
rect 190076 151103 190164 151114
rect 190076 151044 190078 151103
rect 190154 151044 190164 151103
rect 190076 151034 190164 151044
rect 192168 151103 192265 151114
rect 192168 151044 192178 151103
rect 192259 151044 192265 151103
rect 192168 151034 192265 151044
rect 208468 151103 208556 151114
rect 208468 151044 208474 151103
rect 208555 151044 208556 151103
rect 208468 151034 208556 151044
rect 208576 151103 208664 151114
rect 208576 151044 208578 151103
rect 208654 151044 208664 151103
rect 208576 151034 208664 151044
rect 218668 151103 218765 151114
rect 218668 151044 218678 151103
rect 218759 151044 218765 151103
rect 218668 151034 218765 151044
rect 11149 128183 11199 128191
rect 11149 128149 11157 128183
rect 11191 128149 11199 128183
rect 11149 128141 11199 128149
rect 33649 128183 33699 128191
rect 33649 128149 33657 128183
rect 33691 128149 33699 128183
rect 33649 128141 33699 128149
rect 56149 128183 56199 128191
rect 56149 128149 56157 128183
rect 56191 128149 56199 128183
rect 56149 128141 56199 128149
rect 78649 128183 78716 128191
rect 78649 128149 78657 128183
rect 78691 128149 78716 128183
rect 78649 128141 78716 128149
rect 101149 128183 101199 128191
rect 101149 128149 101157 128183
rect 101191 128149 101199 128183
rect 101149 128141 101199 128149
rect 123649 128183 123866 128191
rect 123649 128149 123657 128183
rect 123860 128149 123866 128183
rect 123649 128141 123866 128149
rect 146149 128183 146566 128191
rect 146149 128149 146157 128183
rect 146149 128148 146178 128149
rect 146552 128148 146566 128183
rect 146149 128141 146566 128148
rect 168649 128183 169463 128191
rect 168649 128149 168657 128183
rect 168649 128148 168680 128149
rect 169445 128148 169463 128183
rect 168649 128141 169463 128148
rect 190176 128184 192154 128191
rect 213649 128186 213699 128191
rect 190176 128150 190186 128184
rect 192127 128150 192154 128184
rect 190176 128149 191157 128150
rect 191191 128149 192154 128150
rect 190176 128146 192154 128149
rect 208670 128183 218658 128186
rect 208670 128178 213657 128183
rect 213691 128178 218658 128183
rect 208670 128148 208679 128178
rect 218645 128148 218658 128178
rect 191149 128141 191199 128146
rect 208670 128140 218658 128148
rect 10968 128103 11056 128114
rect 10968 128028 10974 128103
rect 11055 128028 11056 128103
rect 10968 128018 11056 128028
rect 11076 128103 11164 128114
rect 11076 128028 11078 128103
rect 11154 128028 11164 128103
rect 11076 128018 11164 128028
rect 11183 128103 11279 128114
rect 11183 128028 11193 128103
rect 11274 128028 11279 128103
rect 11183 128018 11279 128028
rect 33468 128103 33556 128114
rect 33468 128028 33474 128103
rect 33555 128028 33556 128103
rect 33468 128018 33556 128028
rect 33576 128103 33664 128114
rect 33576 128028 33578 128103
rect 33654 128028 33664 128103
rect 33576 128018 33664 128028
rect 33686 128103 33782 128114
rect 33686 128028 33696 128103
rect 33777 128028 33782 128103
rect 33686 128018 33782 128028
rect 55968 128103 56056 128114
rect 55968 128028 55974 128103
rect 56055 128028 56056 128103
rect 55968 128018 56056 128028
rect 56076 128103 56164 128114
rect 56076 128028 56078 128103
rect 56154 128028 56164 128103
rect 56076 128018 56164 128028
rect 56193 128103 56289 128114
rect 56193 128028 56203 128103
rect 56284 128028 56289 128103
rect 56193 128018 56289 128028
rect 78468 128103 78556 128114
rect 78468 128028 78474 128103
rect 78555 128028 78556 128103
rect 78468 128018 78556 128028
rect 78576 128103 78664 128114
rect 78576 128028 78578 128103
rect 78654 128028 78664 128103
rect 78576 128018 78664 128028
rect 78718 128103 78814 128114
rect 78718 128028 78728 128103
rect 78809 128028 78814 128103
rect 78718 128018 78814 128028
rect 100968 128103 101056 128114
rect 100968 128028 100974 128103
rect 101055 128028 101056 128103
rect 100968 128018 101056 128028
rect 101076 128103 101164 128114
rect 101076 128028 101078 128103
rect 101154 128028 101164 128103
rect 101076 128018 101164 128028
rect 101268 128103 101364 128114
rect 101268 128028 101278 128103
rect 101359 128028 101364 128103
rect 101268 128018 101364 128028
rect 123468 128103 123556 128114
rect 123468 128028 123474 128103
rect 123555 128028 123556 128103
rect 123468 128018 123556 128028
rect 123576 128103 123664 128114
rect 123576 128028 123578 128103
rect 123654 128028 123664 128103
rect 123576 128018 123664 128028
rect 123868 128103 123964 128114
rect 123868 128028 123878 128103
rect 123959 128028 123964 128103
rect 123868 128018 123964 128028
rect 145968 128103 146056 128114
rect 145968 128028 145974 128103
rect 146055 128028 146056 128103
rect 145968 128018 146056 128028
rect 146076 128103 146164 128114
rect 146076 128028 146078 128103
rect 146154 128028 146164 128103
rect 146076 128018 146164 128028
rect 146568 128103 146664 128114
rect 146568 128028 146578 128103
rect 146659 128028 146664 128103
rect 146568 128018 146664 128028
rect 168468 128103 168556 128114
rect 168468 128028 168474 128103
rect 168555 128028 168556 128103
rect 168468 128018 168556 128028
rect 168576 128103 168664 128114
rect 168576 128028 168578 128103
rect 168654 128028 168664 128103
rect 168576 128018 168664 128028
rect 169468 128103 169564 128114
rect 169468 128028 169478 128103
rect 169559 128028 169564 128103
rect 169468 128018 169564 128028
rect 189968 128103 190056 128114
rect 189968 128028 189974 128103
rect 190055 128028 190056 128103
rect 189968 128018 190056 128028
rect 190076 128103 190164 128114
rect 190076 128028 190078 128103
rect 190154 128028 190164 128103
rect 190076 128018 190164 128028
rect 192168 128103 192270 128114
rect 192168 128028 192178 128103
rect 192259 128028 192270 128103
rect 192168 128018 192270 128028
rect 208468 128103 208556 128114
rect 208468 128028 208474 128103
rect 208555 128028 208556 128103
rect 208468 128018 208556 128028
rect 208576 128103 208664 128114
rect 208576 128028 208578 128103
rect 208654 128028 208664 128103
rect 208576 128018 208664 128028
rect 218668 128103 218770 128114
rect 218668 128028 218678 128103
rect 218759 128028 218770 128103
rect 218668 128018 218770 128028
rect 11149 105183 11199 105191
rect 11149 105149 11157 105183
rect 11191 105149 11199 105183
rect 11149 105141 11199 105149
rect 33649 105183 33699 105191
rect 33649 105149 33657 105183
rect 33691 105149 33699 105183
rect 33649 105141 33699 105149
rect 56149 105183 56199 105191
rect 56149 105149 56157 105183
rect 56191 105149 56199 105183
rect 56149 105141 56199 105149
rect 78649 105183 78716 105191
rect 78649 105149 78657 105183
rect 78691 105149 78716 105183
rect 78649 105141 78716 105149
rect 101149 105183 101199 105191
rect 101149 105149 101157 105183
rect 101191 105149 101199 105183
rect 101149 105141 101199 105149
rect 123649 105183 123866 105191
rect 123649 105149 123657 105183
rect 123860 105149 123866 105183
rect 123649 105141 123866 105149
rect 146149 105183 146566 105191
rect 146149 105149 146157 105183
rect 146149 105148 146178 105149
rect 146552 105148 146566 105183
rect 146149 105141 146566 105148
rect 168649 105183 169463 105191
rect 168649 105149 168657 105183
rect 168649 105148 168680 105149
rect 169445 105148 169463 105183
rect 168649 105141 169463 105148
rect 190176 105184 192154 105191
rect 213649 105186 213699 105191
rect 190176 105150 190186 105184
rect 192127 105150 192154 105184
rect 190176 105149 191157 105150
rect 191191 105149 192154 105150
rect 190176 105146 192154 105149
rect 208670 105183 218658 105186
rect 208670 105178 213657 105183
rect 213691 105178 218658 105183
rect 208670 105148 208679 105178
rect 218645 105148 218658 105178
rect 191149 105141 191199 105146
rect 208670 105140 218658 105148
rect 10968 105103 11056 105114
rect 10968 104963 10974 105103
rect 11055 104963 11056 105103
rect 10968 104953 11056 104963
rect 11076 105103 11164 105114
rect 11076 104963 11078 105103
rect 11154 104963 11164 105103
rect 11076 104953 11164 104963
rect 11183 105103 11279 105114
rect 11183 104963 11193 105103
rect 11274 104963 11279 105103
rect 11183 104953 11279 104963
rect 33468 105103 33556 105114
rect 33468 104963 33474 105103
rect 33555 104963 33556 105103
rect 33468 104953 33556 104963
rect 33576 105103 33664 105114
rect 33576 104963 33578 105103
rect 33654 104963 33664 105103
rect 33576 104953 33664 104963
rect 33686 105103 33782 105114
rect 33686 104963 33696 105103
rect 33777 104963 33782 105103
rect 33686 104953 33782 104963
rect 55968 105103 56056 105114
rect 55968 104963 55974 105103
rect 56055 104963 56056 105103
rect 55968 104953 56056 104963
rect 56076 105103 56164 105114
rect 56076 104963 56078 105103
rect 56154 104963 56164 105103
rect 56076 104953 56164 104963
rect 56193 105103 56289 105114
rect 56193 104963 56203 105103
rect 56284 104963 56289 105103
rect 56193 104953 56289 104963
rect 78468 105103 78556 105114
rect 78468 104963 78474 105103
rect 78555 104963 78556 105103
rect 78468 104953 78556 104963
rect 78576 105103 78664 105114
rect 78576 104963 78578 105103
rect 78654 104963 78664 105103
rect 78576 104953 78664 104963
rect 78718 105103 78814 105114
rect 78718 104963 78728 105103
rect 78809 104963 78814 105103
rect 78718 104953 78814 104963
rect 100968 105103 101056 105114
rect 100968 104963 100974 105103
rect 101055 104963 101056 105103
rect 100968 104953 101056 104963
rect 101076 105103 101164 105114
rect 101076 104963 101078 105103
rect 101154 104963 101164 105103
rect 101076 104953 101164 104963
rect 101268 105103 101364 105114
rect 101268 104963 101278 105103
rect 101359 104963 101364 105103
rect 101268 104953 101364 104963
rect 123468 105103 123556 105114
rect 123468 104963 123474 105103
rect 123555 104963 123556 105103
rect 123468 104953 123556 104963
rect 123576 105103 123664 105114
rect 123576 104963 123578 105103
rect 123654 104963 123664 105103
rect 123576 104953 123664 104963
rect 123868 105103 123964 105114
rect 123868 104963 123878 105103
rect 123959 104963 123964 105103
rect 123868 104953 123964 104963
rect 145968 105103 146056 105114
rect 145968 104963 145974 105103
rect 146055 104963 146056 105103
rect 145968 104953 146056 104963
rect 146076 105103 146164 105114
rect 146076 104963 146078 105103
rect 146154 104963 146164 105103
rect 146076 104953 146164 104963
rect 146568 105103 146664 105114
rect 146568 104963 146578 105103
rect 146659 104963 146664 105103
rect 146568 104953 146664 104963
rect 168468 105103 168556 105114
rect 168468 104963 168474 105103
rect 168555 104963 168556 105103
rect 168468 104953 168556 104963
rect 168576 105103 168664 105114
rect 168576 104963 168578 105103
rect 168654 104963 168664 105103
rect 168576 104953 168664 104963
rect 169468 105103 169564 105114
rect 169468 104963 169478 105103
rect 169559 104963 169564 105103
rect 169468 104953 169564 104963
rect 189968 105103 190056 105114
rect 189968 104963 189974 105103
rect 190055 104963 190056 105103
rect 189968 104953 190056 104963
rect 190076 105103 190164 105114
rect 190076 104963 190078 105103
rect 190154 104963 190164 105103
rect 190076 104953 190164 104963
rect 192168 105103 192265 105114
rect 192168 104963 192178 105103
rect 192259 104963 192265 105103
rect 192168 104953 192265 104963
rect 208468 105103 208556 105114
rect 208468 104963 208474 105103
rect 208555 104963 208556 105103
rect 208468 104953 208556 104963
rect 208576 105103 208664 105114
rect 208576 104963 208578 105103
rect 208654 104963 208664 105103
rect 208576 104953 208664 104963
rect 218668 105103 218770 105114
rect 218668 104963 218678 105103
rect 218759 104963 218770 105103
rect 218668 104953 218770 104963
rect 11149 82183 11199 82191
rect 11149 82149 11157 82183
rect 11191 82149 11199 82183
rect 11149 82141 11199 82149
rect 33649 82183 33699 82191
rect 33649 82149 33657 82183
rect 33691 82149 33699 82183
rect 33649 82141 33699 82149
rect 56149 82183 56199 82191
rect 56149 82149 56157 82183
rect 56191 82149 56199 82183
rect 56149 82141 56199 82149
rect 78649 82183 78716 82191
rect 78649 82149 78657 82183
rect 78691 82149 78716 82183
rect 78649 82141 78716 82149
rect 101149 82183 101199 82191
rect 101149 82149 101157 82183
rect 101191 82149 101199 82183
rect 101149 82141 101199 82149
rect 123649 82183 123866 82191
rect 123649 82149 123657 82183
rect 123860 82149 123866 82183
rect 123649 82141 123866 82149
rect 146149 82183 146566 82191
rect 146149 82149 146157 82183
rect 146149 82148 146178 82149
rect 146552 82148 146566 82183
rect 146149 82141 146566 82148
rect 168649 82183 169463 82191
rect 168649 82149 168657 82183
rect 168649 82148 168680 82149
rect 169445 82148 169463 82183
rect 168649 82141 169463 82148
rect 190176 82184 192154 82191
rect 213649 82186 213699 82191
rect 190176 82150 190186 82184
rect 192127 82150 192154 82184
rect 190176 82149 191157 82150
rect 191191 82149 192154 82150
rect 190176 82146 192154 82149
rect 208670 82183 218658 82186
rect 208670 82178 213657 82183
rect 213691 82178 218658 82183
rect 208670 82148 208679 82178
rect 218645 82148 218658 82178
rect 191149 82141 191199 82146
rect 208670 82140 218658 82148
rect 10968 82103 11056 82114
rect 10968 81840 10974 82103
rect 10968 81828 10979 81840
rect 11055 81828 11056 82103
rect 10968 81818 11056 81828
rect 11076 82103 11164 82114
rect 11076 81828 11078 82103
rect 11154 81828 11164 82103
rect 11076 81818 11164 81828
rect 11183 82103 11279 82114
rect 11183 81828 11193 82103
rect 11274 81828 11279 82103
rect 11183 81818 11279 81828
rect 33468 82103 33556 82114
rect 33468 81845 33474 82103
rect 33468 81828 33479 81845
rect 33555 81828 33556 82103
rect 33468 81818 33556 81828
rect 33576 82103 33664 82114
rect 33576 81828 33578 82103
rect 33654 81828 33664 82103
rect 33576 81818 33664 81828
rect 33686 82103 33782 82114
rect 33686 81828 33696 82103
rect 33777 81828 33782 82103
rect 33686 81818 33782 81828
rect 55968 82103 56056 82114
rect 55968 81845 55974 82103
rect 55968 81828 55979 81845
rect 56055 81828 56056 82103
rect 55968 81818 56056 81828
rect 56076 82103 56164 82114
rect 56076 81828 56078 82103
rect 56154 81828 56164 82103
rect 56076 81818 56164 81828
rect 56193 82103 56289 82114
rect 56193 81828 56203 82103
rect 56284 81828 56289 82103
rect 56193 81818 56289 81828
rect 78468 82103 78556 82114
rect 78468 81840 78474 82103
rect 78468 81828 78479 81840
rect 78555 81828 78556 82103
rect 78468 81818 78556 81828
rect 78576 82103 78664 82114
rect 78576 81828 78578 82103
rect 78654 81828 78664 82103
rect 78576 81818 78664 81828
rect 78718 82103 78814 82114
rect 78718 81828 78728 82103
rect 78809 81828 78814 82103
rect 78718 81818 78814 81828
rect 100968 82103 101056 82114
rect 100968 81840 100974 82103
rect 100968 81828 100979 81840
rect 101055 81828 101056 82103
rect 100968 81818 101056 81828
rect 101076 82103 101164 82114
rect 101076 81828 101078 82103
rect 101154 81828 101164 82103
rect 101076 81818 101164 81828
rect 101268 82103 101364 82114
rect 101268 81828 101278 82103
rect 101359 81828 101364 82103
rect 101268 81818 101364 81828
rect 123468 82103 123556 82114
rect 123468 81845 123474 82103
rect 123468 81828 123479 81845
rect 123555 81828 123556 82103
rect 123468 81818 123556 81828
rect 123576 82103 123664 82114
rect 123576 81828 123578 82103
rect 123654 81828 123664 82103
rect 123576 81818 123664 81828
rect 123868 82103 123964 82114
rect 123868 81828 123878 82103
rect 123959 81828 123964 82103
rect 123868 81818 123964 81828
rect 145968 82103 146056 82114
rect 145968 81840 145974 82103
rect 145968 81828 145979 81840
rect 146055 81828 146056 82103
rect 145968 81818 146056 81828
rect 146076 82103 146164 82114
rect 146076 81828 146078 82103
rect 146154 81828 146164 82103
rect 146076 81818 146164 81828
rect 146568 82103 146664 82114
rect 146568 81828 146578 82103
rect 146659 81828 146664 82103
rect 146568 81818 146664 81828
rect 168468 82103 168556 82114
rect 168468 81845 168474 82103
rect 168468 81828 168479 81845
rect 168555 81828 168556 82103
rect 168468 81818 168556 81828
rect 168576 82103 168664 82114
rect 168576 81828 168578 82103
rect 168654 81828 168664 82103
rect 168576 81818 168664 81828
rect 169468 82103 169564 82114
rect 169468 81828 169478 82103
rect 169559 81828 169564 82103
rect 169468 81818 169564 81828
rect 189968 82103 190056 82114
rect 189968 81875 189974 82103
rect 189968 81828 189979 81875
rect 190055 81828 190056 82103
rect 189968 81818 190056 81828
rect 190076 82103 190164 82114
rect 190076 81828 190078 82103
rect 190154 81828 190164 82103
rect 190076 81818 190164 81828
rect 192168 82103 192265 82114
rect 192168 81828 192178 82103
rect 192259 81828 192265 82103
rect 192168 81818 192265 81828
rect 208468 82103 208556 82114
rect 208468 81828 208474 82103
rect 208555 81828 208556 82103
rect 208468 81818 208556 81828
rect 208576 82103 208664 82114
rect 208576 81828 208578 82103
rect 208654 81828 208664 82103
rect 208576 81818 208664 81828
rect 218668 82103 218770 82114
rect 218668 81828 218678 82103
rect 218759 81828 218770 82103
rect 218668 81818 218770 81828
rect 11149 59183 11199 59191
rect 11149 59149 11157 59183
rect 11191 59149 11199 59183
rect 11149 59141 11199 59149
rect 33649 59183 33699 59191
rect 33649 59149 33657 59183
rect 33691 59149 33699 59183
rect 33649 59141 33699 59149
rect 56149 59183 56199 59191
rect 56149 59149 56157 59183
rect 56191 59149 56199 59183
rect 56149 59141 56199 59149
rect 78649 59183 78716 59191
rect 78649 59149 78657 59183
rect 78691 59149 78716 59183
rect 78649 59141 78716 59149
rect 101149 59183 101199 59191
rect 101149 59149 101157 59183
rect 101191 59149 101199 59183
rect 101149 59141 101199 59149
rect 123649 59183 123866 59191
rect 123649 59149 123657 59183
rect 123860 59149 123866 59183
rect 123649 59141 123866 59149
rect 146149 59183 146566 59191
rect 146149 59149 146157 59183
rect 146149 59148 146178 59149
rect 146552 59148 146566 59183
rect 146149 59141 146566 59148
rect 168649 59183 169463 59191
rect 168649 59149 168657 59183
rect 168649 59148 168680 59149
rect 169445 59148 169463 59183
rect 168649 59141 169463 59148
rect 190176 59184 192154 59191
rect 213649 59186 213699 59191
rect 190176 59150 190186 59184
rect 192127 59150 192154 59184
rect 190176 59149 191157 59150
rect 191191 59149 192154 59150
rect 190176 59146 192154 59149
rect 208670 59183 218658 59186
rect 208670 59178 213657 59183
rect 213691 59178 218658 59183
rect 208670 59148 208679 59178
rect 218645 59148 218658 59178
rect 191149 59141 191199 59146
rect 208670 59140 218658 59148
rect 10968 59103 11056 59114
rect 10968 58633 10974 59103
rect 10968 58628 10979 58633
rect 11055 58628 11056 59103
rect 10968 58618 11056 58628
rect 11076 59103 11164 59114
rect 11076 58628 11078 59103
rect 11154 58628 11164 59103
rect 11076 58618 11164 58628
rect 11183 59103 11279 59114
rect 11183 58628 11193 59103
rect 11274 58946 11279 59103
rect 11275 58633 11279 58946
rect 11269 58628 11279 58633
rect 11183 58618 11279 58628
rect 33468 59103 33556 59114
rect 33468 58628 33474 59103
rect 33555 58628 33556 59103
rect 33468 58618 33556 58628
rect 33576 59103 33664 59114
rect 33576 58628 33578 59103
rect 33654 58628 33664 59103
rect 33576 58618 33664 58628
rect 33686 59103 33782 59114
rect 33686 58628 33696 59103
rect 33777 58628 33782 59103
rect 33686 58618 33782 58628
rect 55968 59103 56056 59114
rect 55968 58628 55974 59103
rect 56055 58628 56056 59103
rect 55968 58618 56056 58628
rect 56076 59103 56164 59114
rect 56076 58628 56078 59103
rect 56154 58628 56164 59103
rect 56076 58618 56164 58628
rect 56193 59103 56289 59114
rect 56193 58628 56203 59103
rect 56284 58628 56289 59103
rect 56193 58618 56289 58628
rect 78468 59103 78556 59114
rect 78468 58628 78474 59103
rect 78555 58628 78556 59103
rect 78468 58618 78556 58628
rect 78576 59103 78664 59114
rect 78576 58628 78578 59103
rect 78654 58628 78664 59103
rect 78576 58618 78664 58628
rect 78718 59103 78814 59114
rect 78718 58628 78728 59103
rect 78809 58628 78814 59103
rect 78718 58618 78814 58628
rect 100968 59103 101056 59114
rect 100968 58628 100974 59103
rect 101055 58628 101056 59103
rect 100968 58618 101056 58628
rect 101076 59103 101164 59114
rect 101076 58628 101078 59103
rect 101154 58628 101164 59103
rect 101076 58618 101164 58628
rect 101268 59103 101364 59114
rect 101268 58628 101278 59103
rect 101359 58628 101364 59103
rect 101268 58618 101364 58628
rect 123468 59103 123556 59114
rect 123468 58628 123474 59103
rect 123555 58628 123556 59103
rect 123468 58618 123556 58628
rect 123576 59103 123664 59114
rect 123576 58628 123578 59103
rect 123654 58628 123664 59103
rect 123576 58618 123664 58628
rect 123868 59103 123964 59114
rect 123868 58628 123878 59103
rect 123959 58628 123964 59103
rect 123868 58618 123964 58628
rect 145968 59103 146056 59114
rect 145968 58628 145974 59103
rect 146055 58628 146056 59103
rect 145968 58618 146056 58628
rect 146076 59103 146164 59114
rect 146076 58628 146078 59103
rect 146154 58628 146164 59103
rect 146076 58618 146164 58628
rect 146568 59103 146664 59114
rect 146568 58628 146578 59103
rect 146659 58628 146664 59103
rect 146568 58618 146664 58628
rect 168468 59103 168556 59114
rect 168468 58628 168474 59103
rect 168555 58628 168556 59103
rect 168468 58618 168556 58628
rect 168576 59103 168664 59114
rect 168576 58628 168578 59103
rect 168654 58628 168664 59103
rect 168576 58618 168664 58628
rect 169468 59103 169564 59114
rect 169468 58628 169478 59103
rect 169559 58628 169564 59103
rect 169468 58618 169564 58628
rect 189968 59103 190056 59114
rect 189968 58628 189974 59103
rect 190055 58628 190056 59103
rect 189968 58618 190056 58628
rect 190076 59103 190164 59114
rect 190076 58628 190078 59103
rect 190154 58628 190164 59103
rect 190076 58618 190164 58628
rect 192168 59103 192265 59114
rect 192168 58628 192178 59103
rect 192259 58628 192265 59103
rect 192168 58618 192265 58628
rect 208468 59103 208556 59114
rect 208468 58628 208474 59103
rect 208555 58628 208556 59103
rect 208468 58618 208556 58628
rect 208576 59103 208664 59114
rect 208576 58628 208578 59103
rect 208654 58628 208664 59103
rect 208576 58618 208664 58628
rect 218668 59103 218770 59114
rect 218668 58628 218678 59103
rect 218759 58628 218770 59103
rect 218668 58618 218770 58628
rect 11149 36183 11199 36191
rect 11149 36149 11157 36183
rect 11191 36149 11199 36183
rect 11149 36141 11199 36149
rect 33649 36183 33699 36191
rect 33649 36149 33657 36183
rect 33691 36149 33699 36183
rect 33649 36141 33699 36149
rect 56149 36183 56199 36191
rect 56149 36149 56157 36183
rect 56191 36149 56199 36183
rect 56149 36141 56199 36149
rect 78649 36183 78716 36191
rect 78649 36149 78657 36183
rect 78691 36149 78716 36183
rect 78649 36141 78716 36149
rect 101149 36183 101199 36191
rect 101149 36149 101157 36183
rect 101191 36149 101199 36183
rect 101149 36141 101199 36149
rect 123649 36183 123866 36191
rect 123649 36149 123657 36183
rect 123860 36149 123866 36183
rect 123649 36141 123866 36149
rect 146149 36183 146566 36191
rect 146149 36149 146157 36183
rect 146149 36148 146178 36149
rect 146552 36148 146566 36183
rect 146149 36141 146566 36148
rect 168649 36183 169463 36191
rect 168649 36149 168657 36183
rect 168649 36148 168680 36149
rect 169445 36148 169463 36183
rect 168649 36141 169463 36148
rect 190176 36184 192154 36191
rect 213649 36186 213699 36191
rect 190176 36150 190186 36184
rect 192127 36150 192154 36184
rect 190176 36149 191157 36150
rect 191191 36149 192154 36150
rect 190176 36146 192154 36149
rect 208670 36183 218658 36186
rect 208670 36178 213657 36183
rect 213691 36178 218658 36183
rect 208670 36148 208679 36178
rect 218645 36148 218658 36178
rect 191149 36141 191199 36146
rect 208670 36140 218658 36148
rect 10968 36103 11056 36114
rect 10968 35428 10974 36103
rect 11055 35428 11056 36103
rect 10968 35418 11056 35428
rect 11076 36103 11164 36114
rect 11076 35428 11078 36103
rect 11154 35428 11164 36103
rect 11076 35418 11164 35428
rect 11183 36103 11279 36114
rect 11183 35428 11193 36103
rect 11274 35428 11279 36103
rect 11183 35418 11279 35428
rect 33468 36103 33556 36114
rect 33468 35428 33474 36103
rect 33555 35428 33556 36103
rect 33468 35418 33556 35428
rect 33576 36103 33664 36114
rect 33576 35428 33578 36103
rect 33654 35428 33664 36103
rect 33576 35418 33664 35428
rect 33686 36103 33782 36114
rect 33686 35428 33696 36103
rect 33777 35428 33782 36103
rect 33686 35418 33782 35428
rect 55968 36103 56056 36114
rect 55968 35428 55974 36103
rect 56055 35428 56056 36103
rect 55968 35418 56056 35428
rect 56076 36103 56164 36114
rect 56076 35428 56078 36103
rect 56154 35428 56164 36103
rect 56076 35418 56164 35428
rect 56193 36103 56289 36114
rect 56193 35428 56203 36103
rect 56284 35428 56289 36103
rect 56193 35418 56289 35428
rect 78468 36103 78556 36114
rect 78468 35428 78474 36103
rect 78555 35428 78556 36103
rect 78468 35418 78556 35428
rect 78576 36103 78664 36114
rect 78576 35428 78578 36103
rect 78654 35428 78664 36103
rect 78576 35418 78664 35428
rect 78718 36103 78814 36114
rect 78718 35428 78728 36103
rect 78809 35428 78814 36103
rect 78718 35418 78814 35428
rect 100968 36103 101056 36114
rect 100968 35428 100974 36103
rect 101055 35428 101056 36103
rect 100968 35418 101056 35428
rect 101076 36103 101164 36114
rect 101076 35428 101078 36103
rect 101154 35428 101164 36103
rect 101076 35418 101164 35428
rect 101268 36103 101364 36114
rect 101268 35428 101278 36103
rect 101359 35428 101364 36103
rect 101268 35418 101364 35428
rect 123468 36103 123556 36114
rect 123468 35428 123474 36103
rect 123555 35428 123556 36103
rect 123468 35418 123556 35428
rect 123576 36103 123664 36114
rect 123576 35428 123578 36103
rect 123654 35428 123664 36103
rect 123576 35418 123664 35428
rect 123868 36103 123964 36114
rect 123868 35428 123878 36103
rect 123959 35428 123964 36103
rect 123868 35418 123964 35428
rect 145968 36103 146056 36114
rect 145968 35428 145974 36103
rect 146055 35428 146056 36103
rect 145968 35418 146056 35428
rect 146076 36103 146164 36114
rect 146076 35428 146078 36103
rect 146154 35428 146164 36103
rect 146076 35418 146164 35428
rect 146568 36103 146664 36114
rect 146568 35428 146578 36103
rect 146659 35428 146664 36103
rect 146568 35418 146664 35428
rect 168468 36103 168556 36114
rect 168468 35428 168474 36103
rect 168555 35428 168556 36103
rect 168468 35418 168556 35428
rect 168576 36103 168664 36114
rect 168576 35428 168578 36103
rect 168654 35428 168664 36103
rect 168576 35418 168664 35428
rect 169468 36103 169564 36114
rect 169468 35428 169478 36103
rect 169559 35428 169564 36103
rect 169468 35418 169564 35428
rect 189968 36103 190056 36114
rect 189968 35428 189974 36103
rect 190055 35428 190056 36103
rect 189968 35418 190056 35428
rect 190076 36103 190164 36114
rect 190076 35428 190078 36103
rect 190154 35428 190164 36103
rect 190076 35418 190164 35428
rect 192168 36103 192270 36114
rect 192168 35428 192178 36103
rect 192259 35428 192270 36103
rect 192168 35418 192270 35428
rect 208468 36103 208556 36114
rect 208468 35428 208474 36103
rect 208555 35428 208556 36103
rect 208468 35418 208556 35428
rect 208576 36103 208664 36114
rect 208576 35428 208578 36103
rect 208654 35428 208664 36103
rect 208576 35418 208664 35428
rect 218668 36103 218770 36114
rect 218668 35428 218678 36103
rect 218759 35428 218770 36103
rect 218668 35418 218770 35428
rect 11149 13183 11199 13191
rect 11149 13149 11157 13183
rect 11191 13149 11199 13183
rect 11149 13141 11199 13149
rect 33649 13183 33699 13191
rect 33649 13149 33657 13183
rect 33691 13149 33699 13183
rect 33649 13141 33699 13149
rect 56149 13183 56199 13191
rect 56149 13149 56157 13183
rect 56191 13149 56199 13183
rect 56149 13141 56199 13149
rect 78649 13183 78716 13191
rect 78649 13149 78657 13183
rect 78691 13149 78716 13183
rect 78649 13141 78716 13149
rect 101149 13183 101199 13191
rect 101149 13149 101157 13183
rect 101191 13149 101199 13183
rect 101149 13141 101199 13149
rect 123649 13183 123866 13191
rect 123649 13149 123657 13183
rect 123860 13149 123866 13183
rect 123649 13141 123866 13149
rect 146149 13183 146566 13191
rect 146149 13149 146157 13183
rect 146149 13148 146178 13149
rect 146552 13148 146566 13183
rect 146149 13141 146566 13148
rect 168649 13183 169463 13191
rect 168649 13149 168657 13183
rect 168649 13148 168680 13149
rect 169445 13148 169463 13183
rect 168649 13141 169463 13148
rect 190176 13184 192154 13191
rect 213649 13186 213699 13191
rect 190176 13150 190186 13184
rect 192127 13150 192154 13184
rect 190176 13149 191157 13150
rect 191191 13149 192154 13150
rect 190176 13146 192154 13149
rect 208670 13183 218658 13186
rect 208670 13178 213657 13183
rect 213691 13178 218658 13183
rect 208670 13148 208679 13178
rect 218645 13148 218658 13178
rect 191149 13141 191199 13146
rect 208670 13140 218658 13148
rect 10968 13103 11056 13114
rect 10968 3128 10974 13103
rect 11055 3128 11056 13103
rect 10968 3118 11056 3128
rect 11076 13103 11164 13114
rect 11076 3128 11078 13103
rect 11154 3128 11164 13103
rect 11076 3118 11164 3128
rect 11183 13103 11279 13114
rect 11183 3128 11193 13103
rect 11274 3128 11279 13103
rect 11183 3118 11279 3128
rect 33468 13103 33556 13114
rect 33468 3128 33474 13103
rect 33555 3128 33556 13103
rect 33468 3118 33556 3128
rect 33576 13103 33664 13114
rect 33576 3128 33578 13103
rect 33654 3128 33664 13103
rect 33576 3118 33664 3128
rect 33686 13103 33782 13114
rect 33686 3128 33696 13103
rect 33777 3128 33782 13103
rect 33686 3118 33782 3128
rect 55968 13103 56056 13114
rect 55968 3128 55974 13103
rect 56055 3128 56056 13103
rect 55968 3118 56056 3128
rect 56076 13103 56164 13114
rect 56076 3128 56078 13103
rect 56154 3128 56164 13103
rect 56076 3118 56164 3128
rect 56193 13103 56289 13114
rect 56193 3128 56203 13103
rect 56284 3128 56289 13103
rect 56193 3118 56289 3128
rect 78468 13103 78556 13114
rect 78468 3128 78474 13103
rect 78555 3128 78556 13103
rect 78468 3118 78556 3128
rect 78576 13103 78664 13114
rect 78576 3128 78578 13103
rect 78654 3128 78664 13103
rect 78576 3118 78664 3128
rect 78718 13103 78814 13114
rect 78718 3128 78728 13103
rect 78809 3128 78814 13103
rect 78718 3118 78814 3128
rect 100968 13103 101056 13114
rect 100968 3128 100974 13103
rect 101055 3128 101056 13103
rect 100968 3118 101056 3128
rect 101076 13103 101164 13114
rect 101076 3128 101078 13103
rect 101154 3128 101164 13103
rect 101076 3118 101164 3128
rect 101268 13103 101364 13114
rect 101268 3128 101278 13103
rect 101359 3128 101364 13103
rect 101268 3118 101364 3128
rect 123468 13103 123556 13114
rect 123468 3128 123474 13103
rect 123555 3128 123556 13103
rect 123468 3118 123556 3128
rect 123576 13103 123664 13114
rect 123576 3128 123578 13103
rect 123654 3128 123664 13103
rect 123576 3118 123664 3128
rect 123868 13103 123964 13114
rect 123868 3128 123878 13103
rect 123959 3128 123964 13103
rect 123868 3118 123964 3128
rect 145968 13103 146056 13114
rect 145968 3128 145974 13103
rect 146055 3128 146056 13103
rect 145968 3118 146056 3128
rect 146076 13103 146164 13114
rect 146076 3128 146078 13103
rect 146154 3128 146164 13103
rect 146076 3118 146164 3128
rect 146568 13103 146664 13114
rect 146568 3128 146578 13103
rect 146659 3128 146664 13103
rect 146568 3118 146664 3128
rect 168468 13103 168556 13114
rect 168468 3128 168474 13103
rect 168555 3128 168556 13103
rect 168468 3118 168556 3128
rect 168576 13103 168664 13114
rect 168576 3128 168578 13103
rect 168654 3128 168664 13103
rect 168576 3118 168664 3128
rect 169468 13103 169564 13114
rect 169468 3128 169478 13103
rect 169559 3128 169564 13103
rect 169468 3118 169564 3128
rect 189968 13103 190056 13114
rect 189968 3128 189974 13103
rect 190055 3128 190056 13103
rect 189968 3118 190056 3128
rect 190076 13103 190164 13114
rect 190076 3128 190078 13103
rect 190154 3128 190164 13103
rect 190076 3118 190164 3128
rect 192168 13103 192270 13114
rect 192168 3128 192178 13103
rect 192259 3128 192270 13103
rect 192168 3118 192270 3128
rect 208468 13103 208556 13114
rect 208468 3128 208474 13103
rect 208555 3128 208556 13103
rect 208468 3118 208556 3128
rect 208576 13103 208664 13114
rect 208576 3128 208578 13103
rect 208654 3128 208664 13103
rect 208576 3118 208664 3128
rect 218668 13103 218770 13114
rect 218668 3128 218678 13103
rect 218759 3128 218770 13103
rect 218668 3118 218770 3128
<< viali >>
rect 11157 220150 11191 220183
rect 33657 220150 33691 220183
rect 56157 220150 56191 220183
rect 78657 220150 78691 220183
rect 101157 220150 101191 220183
rect 123657 220150 123860 220183
rect 123691 220149 123860 220150
rect 146157 220150 146552 220183
rect 146178 220148 146552 220150
rect 168657 220150 169445 220183
rect 168680 220148 169445 220150
rect 190186 220150 192127 220184
rect 213657 220178 213691 220183
rect 208679 220148 218645 220178
rect 10974 220086 10979 220103
rect 10979 220086 11038 220103
rect 11083 220086 11147 220103
rect 11199 220086 11269 220103
rect 11269 220086 11274 220103
rect 33474 220086 33479 220103
rect 33479 220086 33538 220103
rect 33583 220086 33647 220103
rect 33702 220086 33772 220103
rect 33772 220086 33777 220103
rect 55974 220086 55979 220103
rect 55979 220086 56038 220103
rect 56083 220086 56147 220103
rect 56209 220086 56279 220103
rect 56279 220086 56284 220103
rect 78474 220086 78479 220103
rect 78479 220086 78538 220103
rect 78583 220086 78647 220103
rect 78734 220086 78804 220103
rect 78804 220086 78809 220103
rect 100974 220086 100979 220103
rect 100979 220086 101038 220103
rect 101083 220086 101147 220103
rect 101284 220086 101354 220103
rect 101354 220086 101359 220103
rect 123474 220086 123479 220103
rect 123479 220086 123538 220103
rect 123583 220086 123647 220103
rect 123884 220086 123954 220103
rect 123954 220086 123959 220103
rect 145974 220086 145979 220103
rect 145979 220086 146038 220103
rect 146083 220086 146147 220103
rect 146584 220086 146654 220103
rect 146654 220086 146659 220103
rect 168474 220086 168479 220103
rect 168479 220086 168538 220103
rect 168583 220086 168647 220103
rect 169484 220086 169554 220103
rect 169554 220086 169559 220103
rect 189974 220086 189979 220103
rect 189979 220086 190038 220103
rect 190083 220086 190147 220103
rect 192184 220086 192254 220103
rect 192254 220086 192259 220103
rect 208474 220086 208479 220103
rect 208479 220086 208538 220103
rect 208583 220086 208647 220103
rect 218684 220086 218754 220103
rect 218754 220086 218759 220103
rect 11157 197150 11191 197183
rect 33657 197150 33691 197183
rect 56157 197150 56191 197183
rect 78657 197150 78691 197183
rect 101157 197150 101191 197183
rect 123657 197150 123860 197183
rect 123691 197149 123860 197150
rect 146157 197150 146552 197183
rect 146178 197148 146552 197150
rect 168657 197150 169445 197183
rect 168680 197148 169445 197150
rect 190186 197150 192127 197184
rect 213657 197178 213691 197183
rect 208679 197148 218645 197178
rect 10974 197073 10979 197103
rect 10979 197073 11038 197103
rect 11083 197073 11147 197103
rect 11199 197073 11269 197103
rect 11269 197073 11274 197103
rect 33474 197073 33479 197103
rect 33479 197073 33538 197103
rect 33583 197073 33647 197103
rect 33702 197073 33772 197103
rect 33772 197073 33777 197103
rect 55974 197073 55979 197103
rect 55979 197073 56038 197103
rect 56083 197073 56147 197103
rect 56209 197073 56279 197103
rect 56279 197073 56284 197103
rect 78474 197073 78479 197103
rect 78479 197073 78538 197103
rect 78583 197073 78647 197103
rect 78734 197073 78804 197103
rect 78804 197073 78809 197103
rect 100974 197073 100979 197103
rect 100979 197073 101038 197103
rect 101083 197073 101147 197103
rect 101284 197073 101354 197103
rect 101354 197073 101359 197103
rect 123474 197073 123479 197103
rect 123479 197073 123538 197103
rect 123583 197073 123647 197103
rect 123884 197073 123954 197103
rect 123954 197073 123959 197103
rect 145974 197073 145979 197103
rect 145979 197073 146038 197103
rect 146083 197073 146147 197103
rect 146584 197073 146654 197103
rect 146654 197073 146659 197103
rect 168474 197073 168479 197103
rect 168479 197073 168538 197103
rect 168583 197073 168647 197103
rect 169484 197073 169554 197103
rect 169554 197073 169559 197103
rect 189974 197073 189979 197103
rect 189979 197073 190038 197103
rect 190083 197073 190147 197103
rect 192184 197073 192254 197103
rect 192254 197073 192259 197103
rect 208474 197073 208479 197103
rect 208479 197073 208538 197103
rect 208583 197073 208647 197103
rect 218684 197073 218754 197103
rect 218754 197073 218759 197103
rect 11157 174150 11191 174183
rect 33657 174150 33691 174183
rect 56157 174150 56191 174183
rect 78657 174150 78691 174183
rect 101157 174150 101191 174183
rect 123657 174150 123860 174183
rect 123691 174149 123860 174150
rect 146157 174150 146552 174183
rect 146178 174148 146552 174150
rect 168657 174150 169445 174183
rect 168680 174148 169445 174150
rect 190186 174150 192127 174184
rect 213657 174178 213691 174183
rect 208679 174148 218645 174178
rect 10974 174064 10979 174103
rect 10979 174064 11038 174103
rect 11083 174064 11147 174103
rect 11199 174064 11269 174103
rect 11269 174064 11274 174103
rect 33474 174064 33479 174103
rect 33479 174064 33538 174103
rect 33583 174064 33647 174103
rect 33702 174064 33772 174103
rect 33772 174064 33777 174103
rect 55974 174064 55979 174103
rect 55979 174064 56038 174103
rect 56083 174064 56147 174103
rect 56209 174064 56279 174103
rect 56279 174064 56284 174103
rect 78474 174064 78479 174103
rect 78479 174064 78538 174103
rect 78583 174064 78647 174103
rect 78734 174064 78804 174103
rect 78804 174064 78809 174103
rect 100974 174064 100979 174103
rect 100979 174064 101038 174103
rect 101083 174064 101147 174103
rect 101284 174064 101354 174103
rect 101354 174064 101359 174103
rect 123474 174064 123479 174103
rect 123479 174064 123538 174103
rect 123583 174064 123647 174103
rect 123884 174064 123954 174103
rect 123954 174064 123959 174103
rect 145974 174064 145979 174103
rect 145979 174064 146038 174103
rect 146083 174064 146147 174103
rect 146584 174064 146654 174103
rect 146654 174064 146659 174103
rect 168474 174064 168479 174103
rect 168479 174064 168538 174103
rect 168583 174064 168647 174103
rect 169484 174064 169554 174103
rect 169554 174064 169559 174103
rect 189974 174064 189979 174103
rect 189979 174064 190038 174103
rect 190083 174064 190147 174103
rect 192184 174064 192254 174103
rect 192254 174064 192259 174103
rect 208474 174064 208479 174103
rect 208479 174064 208538 174103
rect 208583 174064 208647 174103
rect 218684 174064 218754 174103
rect 218754 174064 218759 174103
rect 11157 151150 11191 151183
rect 33657 151150 33691 151183
rect 56157 151150 56191 151183
rect 78657 151150 78691 151183
rect 101157 151150 101191 151183
rect 123657 151150 123860 151183
rect 123691 151149 123860 151150
rect 146157 151150 146552 151183
rect 146178 151148 146552 151150
rect 168657 151150 169445 151183
rect 168680 151148 169445 151150
rect 190186 151150 192127 151184
rect 213657 151178 213691 151183
rect 208679 151148 218645 151178
rect 10974 151044 10979 151103
rect 10979 151044 11038 151103
rect 11083 151044 11147 151103
rect 11199 151044 11269 151103
rect 11269 151044 11274 151103
rect 33474 151044 33479 151103
rect 33479 151044 33538 151103
rect 33583 151044 33647 151103
rect 33702 151044 33772 151103
rect 33772 151044 33777 151103
rect 55974 151044 55979 151103
rect 55979 151044 56038 151103
rect 56083 151044 56147 151103
rect 56209 151044 56279 151103
rect 56279 151044 56284 151103
rect 78474 151044 78479 151103
rect 78479 151044 78538 151103
rect 78583 151044 78647 151103
rect 78734 151044 78804 151103
rect 78804 151044 78809 151103
rect 100974 151044 100979 151103
rect 100979 151044 101038 151103
rect 101083 151044 101147 151103
rect 101284 151044 101354 151103
rect 101354 151044 101359 151103
rect 123474 151044 123479 151103
rect 123479 151044 123538 151103
rect 123583 151044 123647 151103
rect 123884 151044 123954 151103
rect 123954 151044 123959 151103
rect 145974 151044 145979 151103
rect 145979 151044 146038 151103
rect 146083 151044 146147 151103
rect 146584 151044 146654 151103
rect 146654 151044 146659 151103
rect 168474 151044 168479 151103
rect 168479 151044 168538 151103
rect 168583 151044 168647 151103
rect 169484 151044 169554 151103
rect 169554 151044 169559 151103
rect 189974 151044 189979 151103
rect 189979 151044 190038 151103
rect 190083 151044 190147 151103
rect 192184 151044 192254 151103
rect 192254 151044 192259 151103
rect 208474 151044 208479 151103
rect 208479 151044 208538 151103
rect 208583 151044 208647 151103
rect 218684 151044 218754 151103
rect 218754 151044 218759 151103
rect 11157 128150 11191 128183
rect 33657 128150 33691 128183
rect 56157 128150 56191 128183
rect 78657 128150 78691 128183
rect 101157 128150 101191 128183
rect 123657 128150 123860 128183
rect 123691 128149 123860 128150
rect 146157 128150 146552 128183
rect 146178 128148 146552 128150
rect 168657 128150 169445 128183
rect 168680 128148 169445 128150
rect 190186 128150 192127 128184
rect 213657 128178 213691 128183
rect 208679 128148 218645 128178
rect 10974 128028 10979 128103
rect 10979 128028 11038 128103
rect 11083 128028 11147 128103
rect 11199 128028 11269 128103
rect 11269 128028 11274 128103
rect 33474 128028 33479 128103
rect 33479 128028 33538 128103
rect 33583 128028 33647 128103
rect 33702 128028 33772 128103
rect 33772 128028 33777 128103
rect 55974 128028 55979 128103
rect 55979 128028 56038 128103
rect 56083 128028 56147 128103
rect 56209 128028 56279 128103
rect 56279 128028 56284 128103
rect 78474 128028 78479 128103
rect 78479 128028 78538 128103
rect 78583 128028 78647 128103
rect 78734 128028 78804 128103
rect 78804 128028 78809 128103
rect 100974 128028 100979 128103
rect 100979 128028 101038 128103
rect 101083 128028 101147 128103
rect 101284 128028 101354 128103
rect 101354 128028 101359 128103
rect 123474 128028 123479 128103
rect 123479 128028 123538 128103
rect 123583 128028 123647 128103
rect 123884 128028 123954 128103
rect 123954 128028 123959 128103
rect 145974 128028 145979 128103
rect 145979 128028 146038 128103
rect 146083 128028 146147 128103
rect 146584 128028 146654 128103
rect 146654 128028 146659 128103
rect 168474 128028 168479 128103
rect 168479 128028 168538 128103
rect 168583 128028 168647 128103
rect 169484 128028 169554 128103
rect 169554 128028 169559 128103
rect 189974 128028 189979 128103
rect 189979 128028 190038 128103
rect 190083 128028 190147 128103
rect 192184 128028 192254 128103
rect 192254 128028 192259 128103
rect 208474 128028 208479 128103
rect 208479 128028 208538 128103
rect 208583 128028 208647 128103
rect 218684 128028 218754 128103
rect 218754 128028 218759 128103
rect 11157 105150 11191 105183
rect 33657 105150 33691 105183
rect 56157 105150 56191 105183
rect 78657 105150 78691 105183
rect 101157 105150 101191 105183
rect 123657 105150 123860 105183
rect 123691 105149 123860 105150
rect 146157 105150 146552 105183
rect 146178 105148 146552 105150
rect 168657 105150 169445 105183
rect 168680 105148 169445 105150
rect 190186 105150 192127 105184
rect 213657 105178 213691 105183
rect 208679 105148 218645 105178
rect 10974 104963 10979 105103
rect 10979 104963 11038 105103
rect 11083 104963 11147 105103
rect 11199 104963 11269 105103
rect 11269 104963 11274 105103
rect 33474 104963 33479 105103
rect 33479 104963 33538 105103
rect 33583 104963 33647 105103
rect 33702 104963 33772 105103
rect 33772 104963 33777 105103
rect 55974 104963 55979 105103
rect 55979 104963 56038 105103
rect 56083 104963 56147 105103
rect 56209 104963 56279 105103
rect 56279 104963 56284 105103
rect 78474 104963 78479 105103
rect 78479 104963 78538 105103
rect 78583 104963 78647 105103
rect 78734 104963 78804 105103
rect 78804 104963 78809 105103
rect 100974 104963 100979 105103
rect 100979 104963 101038 105103
rect 101083 104963 101147 105103
rect 101284 104963 101354 105103
rect 101354 104963 101359 105103
rect 123474 104963 123479 105103
rect 123479 104963 123538 105103
rect 123583 104963 123647 105103
rect 123884 104963 123954 105103
rect 123954 104963 123959 105103
rect 145974 104963 145979 105103
rect 145979 104963 146038 105103
rect 146083 104963 146147 105103
rect 146584 104963 146654 105103
rect 146654 104963 146659 105103
rect 168474 104963 168479 105103
rect 168479 104963 168538 105103
rect 168583 104963 168647 105103
rect 169484 104963 169554 105103
rect 169554 104963 169559 105103
rect 189974 104963 189979 105103
rect 189979 104963 190038 105103
rect 190083 104963 190147 105103
rect 192184 104963 192254 105103
rect 192254 104963 192259 105103
rect 208474 104963 208479 105103
rect 208479 104963 208538 105103
rect 208583 104963 208647 105103
rect 218684 104963 218754 105103
rect 218754 104963 218759 105103
rect 11157 82150 11191 82183
rect 33657 82150 33691 82183
rect 56157 82150 56191 82183
rect 78657 82150 78691 82183
rect 101157 82150 101191 82183
rect 123657 82150 123860 82183
rect 123691 82149 123860 82150
rect 146157 82150 146552 82183
rect 146178 82148 146552 82150
rect 168657 82150 169445 82183
rect 168680 82148 169445 82150
rect 190186 82150 192127 82184
rect 213657 82178 213691 82183
rect 208679 82148 218645 82178
rect 10974 81840 10979 82103
rect 10979 81840 11038 82103
rect 11083 81828 11147 82103
rect 11199 81828 11269 82103
rect 11269 81828 11274 82103
rect 33474 81845 33479 82103
rect 33479 81845 33538 82103
rect 33583 81828 33647 82103
rect 33702 81828 33772 82103
rect 33772 81828 33777 82103
rect 55974 81845 55979 82103
rect 55979 81845 56038 82103
rect 56083 81828 56147 82103
rect 56209 81828 56279 82103
rect 56279 81828 56284 82103
rect 78474 81840 78479 82103
rect 78479 81840 78538 82103
rect 78583 81828 78647 82103
rect 78734 81828 78804 82103
rect 78804 81828 78809 82103
rect 100974 81840 100979 82103
rect 100979 81840 101038 82103
rect 101083 81828 101147 82103
rect 101284 81828 101354 82103
rect 101354 81828 101359 82103
rect 123474 81845 123479 82103
rect 123479 81845 123538 82103
rect 123583 81828 123647 82103
rect 123884 81828 123954 82103
rect 123954 81828 123959 82103
rect 145974 81840 145979 82103
rect 145979 81840 146038 82103
rect 146083 81828 146147 82103
rect 146584 81828 146654 82103
rect 146654 81828 146659 82103
rect 168474 81845 168479 82103
rect 168479 81845 168538 82103
rect 168583 81828 168647 82103
rect 169484 81828 169554 82103
rect 169554 81828 169559 82103
rect 189974 81875 189979 82103
rect 189979 81875 190038 82103
rect 190083 81828 190147 82103
rect 192184 81828 192254 82103
rect 192254 81828 192259 82103
rect 208474 81828 208479 82103
rect 208479 81828 208538 82103
rect 208583 81828 208647 82103
rect 218684 81828 218754 82103
rect 218754 81828 218759 82103
rect 11157 59150 11191 59183
rect 33657 59150 33691 59183
rect 56157 59150 56191 59183
rect 78657 59150 78691 59183
rect 101157 59150 101191 59183
rect 123657 59150 123860 59183
rect 123691 59149 123860 59150
rect 146157 59150 146552 59183
rect 146178 59148 146552 59150
rect 168657 59150 169445 59183
rect 168680 59148 169445 59150
rect 190186 59150 192127 59184
rect 213657 59178 213691 59183
rect 208679 59148 218645 59178
rect 10974 58943 10979 59103
rect 10979 58943 11038 59103
rect 10974 58633 11039 58943
rect 11083 58943 11147 59103
rect 11083 58633 11148 58943
rect 11199 58946 11269 59103
rect 11269 58946 11274 59103
rect 11199 58633 11275 58946
rect 33474 58628 33479 59103
rect 33479 58628 33538 59103
rect 33583 58628 33647 59103
rect 33702 58628 33772 59103
rect 33772 58628 33777 59103
rect 55974 58628 55979 59103
rect 55979 58628 56038 59103
rect 56083 58628 56147 59103
rect 56209 58628 56279 59103
rect 56279 58628 56284 59103
rect 78474 58628 78479 59103
rect 78479 58628 78538 59103
rect 78583 58628 78647 59103
rect 78734 58628 78804 59103
rect 78804 58628 78809 59103
rect 100974 58628 100979 59103
rect 100979 58628 101038 59103
rect 101083 58628 101147 59103
rect 101284 58628 101354 59103
rect 101354 58628 101359 59103
rect 123474 58628 123479 59103
rect 123479 58628 123538 59103
rect 123583 58628 123647 59103
rect 123884 58628 123954 59103
rect 123954 58628 123959 59103
rect 145974 58628 145979 59103
rect 145979 58628 146038 59103
rect 146083 58628 146147 59103
rect 146584 58628 146654 59103
rect 146654 58628 146659 59103
rect 168474 58628 168479 59103
rect 168479 58628 168538 59103
rect 168583 58628 168647 59103
rect 169484 58628 169554 59103
rect 169554 58628 169559 59103
rect 189974 58628 189979 59103
rect 189979 58628 190038 59103
rect 190083 58628 190147 59103
rect 192184 58628 192254 59103
rect 192254 58628 192259 59103
rect 208474 58628 208479 59103
rect 208479 58628 208538 59103
rect 208583 58628 208647 59103
rect 218684 58628 218754 59103
rect 218754 58628 218759 59103
rect 11157 36150 11191 36183
rect 33657 36150 33691 36183
rect 56157 36150 56191 36183
rect 78657 36150 78691 36183
rect 101157 36150 101191 36183
rect 123657 36150 123860 36183
rect 123691 36149 123860 36150
rect 146157 36150 146552 36183
rect 146178 36148 146552 36150
rect 168657 36150 169445 36183
rect 168680 36148 169445 36150
rect 190186 36150 192127 36184
rect 213657 36178 213691 36183
rect 208679 36148 218645 36178
rect 10974 35428 10979 36103
rect 10979 35428 11038 36103
rect 11083 35428 11147 36103
rect 11199 35428 11269 36103
rect 11269 35428 11274 36103
rect 33474 35428 33479 36103
rect 33479 35428 33538 36103
rect 33583 35428 33647 36103
rect 33702 35428 33772 36103
rect 33772 35428 33777 36103
rect 55974 35428 55979 36103
rect 55979 35428 56038 36103
rect 56083 35428 56147 36103
rect 56209 35428 56279 36103
rect 56279 35428 56284 36103
rect 78474 35428 78479 36103
rect 78479 35428 78538 36103
rect 78583 35428 78647 36103
rect 78734 35428 78804 36103
rect 78804 35428 78809 36103
rect 100974 35428 100979 36103
rect 100979 35428 101038 36103
rect 101083 35428 101147 36103
rect 101284 35428 101354 36103
rect 101354 35428 101359 36103
rect 123474 35428 123479 36103
rect 123479 35428 123538 36103
rect 123583 35428 123647 36103
rect 123884 35428 123954 36103
rect 123954 35428 123959 36103
rect 145974 35428 145979 36103
rect 145979 35428 146038 36103
rect 146083 35428 146147 36103
rect 146584 35428 146654 36103
rect 146654 35428 146659 36103
rect 168474 35428 168479 36103
rect 168479 35428 168538 36103
rect 168583 35428 168647 36103
rect 169484 35428 169554 36103
rect 169554 35428 169559 36103
rect 189974 35428 189979 36103
rect 189979 35428 190038 36103
rect 190083 35428 190147 36103
rect 192184 35428 192254 36103
rect 192254 35428 192259 36103
rect 208474 35428 208479 36103
rect 208479 35428 208538 36103
rect 208583 35428 208647 36103
rect 218684 35428 218754 36103
rect 218754 35428 218759 36103
rect 11157 13150 11191 13183
rect 33657 13150 33691 13183
rect 56157 13150 56191 13183
rect 78657 13150 78691 13183
rect 101157 13150 101191 13183
rect 123657 13150 123860 13183
rect 123691 13149 123860 13150
rect 146157 13150 146552 13183
rect 146178 13148 146552 13150
rect 168657 13150 169445 13183
rect 168680 13148 169445 13150
rect 190186 13150 192127 13184
rect 213657 13178 213691 13183
rect 208679 13148 218645 13178
rect 10974 3128 10979 13103
rect 10979 3128 11038 13103
rect 11083 3128 11147 13103
rect 11199 3128 11269 13103
rect 11269 3128 11274 13103
rect 33474 3128 33479 13103
rect 33479 3128 33538 13103
rect 33583 3128 33647 13103
rect 33702 3128 33772 13103
rect 33772 3128 33777 13103
rect 55974 3128 55979 13103
rect 55979 3128 56038 13103
rect 56083 3128 56147 13103
rect 56209 3128 56279 13103
rect 56279 3128 56284 13103
rect 78474 3128 78479 13103
rect 78479 3128 78538 13103
rect 78583 3128 78647 13103
rect 78734 3128 78804 13103
rect 78804 3128 78809 13103
rect 100974 3128 100979 13103
rect 100979 3128 101038 13103
rect 101083 3128 101147 13103
rect 101284 3128 101354 13103
rect 101354 3128 101359 13103
rect 123474 3128 123479 13103
rect 123479 3128 123538 13103
rect 123583 3128 123647 13103
rect 123884 3128 123954 13103
rect 123954 3128 123959 13103
rect 145974 3128 145979 13103
rect 145979 3128 146038 13103
rect 146083 3128 146147 13103
rect 146584 3128 146654 13103
rect 146654 3128 146659 13103
rect 168474 3128 168479 13103
rect 168479 3128 168538 13103
rect 168583 3128 168647 13103
rect 169484 3128 169554 13103
rect 169554 3128 169559 13103
rect 189974 3128 189979 13103
rect 189979 3128 190038 13103
rect 190083 3128 190147 13103
rect 192184 3128 192254 13103
rect 192254 3128 192259 13103
rect 208474 3128 208479 13103
rect 208479 3128 208538 13103
rect 208583 3128 208647 13103
rect 218684 3128 218754 13103
rect 218754 3128 218759 13103
<< metal1 >>
rect 10792 220560 11045 221020
rect 10968 220307 11045 220560
rect 32245 220515 33745 221020
rect 54745 220515 56245 221020
rect 77245 220515 78745 221020
rect 99745 220515 101245 221020
rect 122245 220515 123745 221020
rect 144745 220515 146245 221020
rect 167245 220515 168745 221020
rect 189745 220736 191245 221020
rect 189745 220515 190941 220736
rect 191091 220515 191245 220736
rect 33468 220307 33545 220515
rect 55968 220307 56045 220515
rect 78468 220307 78545 220515
rect 100968 220307 101045 220515
rect 123468 220307 123545 220515
rect 145968 220307 146045 220515
rect 168468 220307 168545 220515
rect 10968 220103 11046 220307
rect 11149 220183 13100 220203
rect 11149 220150 11157 220183
rect 11191 220150 13100 220183
rect 11149 220141 13100 220150
rect 10968 220086 10974 220103
rect 11038 220086 11046 220103
rect 10968 220077 11046 220086
rect 11076 220103 11154 220113
rect 11076 220086 11083 220103
rect 11147 220086 11154 220103
rect 11076 219916 11154 220086
rect 11075 219896 11154 219916
rect 11193 220103 11281 220114
rect 11193 220086 11199 220103
rect 11274 220086 11281 220103
rect 11193 220071 11281 220086
rect 33468 220103 33546 220307
rect 33649 220183 35519 220203
rect 33649 220150 33657 220183
rect 33691 220150 35519 220183
rect 33649 220141 35519 220150
rect 33468 220086 33474 220103
rect 33538 220086 33546 220103
rect 33468 220077 33546 220086
rect 33576 220103 33654 220113
rect 33576 220086 33583 220103
rect 33647 220086 33654 220103
rect 11075 219839 11153 219896
rect 10873 219771 11153 219839
rect 11193 219853 11271 220071
rect 33576 219916 33654 220086
rect 33696 220103 33784 220114
rect 33696 220086 33702 220103
rect 33777 220086 33784 220103
rect 33696 220071 33784 220086
rect 55968 220103 56046 220307
rect 57750 220203 58024 220204
rect 56149 220183 58024 220203
rect 56149 220150 56157 220183
rect 56191 220150 58024 220183
rect 56149 220141 58024 220150
rect 55968 220086 55974 220103
rect 56038 220086 56046 220103
rect 55968 220077 56046 220086
rect 56076 220103 56154 220113
rect 56076 220086 56083 220103
rect 56147 220086 56154 220103
rect 33696 220059 33774 220071
rect 33696 220018 33771 220059
rect 33575 219896 33654 219916
rect 11193 219802 11691 219853
rect 33575 219839 33653 219896
rect 10873 219763 11152 219771
rect 10208 219762 11152 219763
rect 8981 219728 11152 219762
rect 11194 219733 11691 219802
rect 33373 219771 33653 219839
rect 33693 219853 33771 220018
rect 56076 219916 56154 220086
rect 56075 219896 56154 219916
rect 56203 220103 56291 220114
rect 56203 220086 56209 220103
rect 56284 220086 56291 220103
rect 56203 220071 56291 220086
rect 78468 220103 78546 220307
rect 78649 220183 80532 220203
rect 78649 220150 78657 220183
rect 78691 220150 80532 220183
rect 78649 220141 80532 220150
rect 78468 220086 78474 220103
rect 78538 220086 78546 220103
rect 78468 220077 78546 220086
rect 78576 220103 78654 220113
rect 78576 220086 78583 220103
rect 78647 220086 78654 220103
rect 33693 219802 34191 219853
rect 56075 219839 56153 219896
rect 8981 219504 10949 219728
rect 11074 219725 11152 219728
rect 8980 219321 10949 219504
rect 8980 219319 10224 219321
rect 8980 218108 9482 219319
rect 11256 215985 11691 219733
rect 31479 219762 32255 219764
rect 33373 219763 33652 219771
rect 32708 219762 33652 219763
rect 31479 219728 33652 219762
rect 33694 219733 34191 219802
rect 55873 219771 56153 219839
rect 56203 219853 56281 220071
rect 78576 219916 78654 220086
rect 78575 219896 78654 219916
rect 78728 220103 78816 220114
rect 78728 220086 78734 220103
rect 78809 220086 78816 220103
rect 78728 220071 78816 220086
rect 100968 220103 101046 220307
rect 101149 220183 103018 220203
rect 101149 220150 101157 220183
rect 101191 220150 103018 220183
rect 101149 220141 103018 220150
rect 100968 220086 100974 220103
rect 101038 220086 101046 220103
rect 100968 220077 101046 220086
rect 101076 220103 101154 220113
rect 101076 220086 101083 220103
rect 101147 220086 101154 220103
rect 56203 219802 56691 219853
rect 78575 219839 78653 219896
rect 55873 219763 56152 219771
rect 55208 219762 56152 219763
rect 31479 219321 33449 219728
rect 33574 219725 33652 219728
rect 31479 219319 32724 219321
rect 31479 218249 32255 219319
rect 33756 216632 34191 219733
rect 53983 219755 54481 219761
rect 54745 219755 56152 219762
rect 53983 219728 56152 219755
rect 56204 219733 56691 219802
rect 78373 219771 78653 219839
rect 78728 219853 78806 220071
rect 101076 219916 101154 220086
rect 101278 220103 101366 220114
rect 101278 220086 101284 220103
rect 101359 220086 101366 220103
rect 101278 220071 101366 220086
rect 123468 220103 123546 220307
rect 123649 220183 125532 220203
rect 123649 220150 123657 220183
rect 123649 220149 123691 220150
rect 123860 220149 125532 220183
rect 123649 220141 125532 220149
rect 125242 220140 125532 220141
rect 123468 220086 123474 220103
rect 123538 220086 123546 220103
rect 123468 220077 123546 220086
rect 123576 220103 123654 220113
rect 123576 220086 123583 220103
rect 123647 220086 123654 220103
rect 101278 220031 101356 220071
rect 101075 219896 101154 219916
rect 78728 219802 79191 219853
rect 101075 219839 101153 219896
rect 101277 219853 101357 220031
rect 123576 219916 123654 220086
rect 123575 219896 123654 219916
rect 123878 220103 123966 220114
rect 123878 220086 123884 220103
rect 123959 220098 123966 220103
rect 145968 220103 146046 220307
rect 146149 220183 148021 220203
rect 146149 220150 146157 220183
rect 146149 220148 146178 220150
rect 146552 220148 148021 220183
rect 146149 220141 148021 220148
rect 123959 220086 123971 220098
rect 53983 219327 55949 219728
rect 56074 219725 56152 219728
rect 56225 219626 56691 219733
rect 53983 218185 54481 219327
rect 54745 219321 55949 219327
rect 54745 219319 55224 219321
rect 56256 216767 56691 219626
rect 76480 219761 76989 219764
rect 78373 219763 78652 219771
rect 77708 219762 78652 219763
rect 77245 219761 78652 219762
rect 76480 219728 78652 219761
rect 78729 219733 79191 219802
rect 100873 219771 101153 219839
rect 100873 219763 101152 219771
rect 100208 219762 101152 219763
rect 99745 219760 101152 219762
rect 99230 219750 101152 219760
rect 76480 219321 78449 219728
rect 78574 219725 78652 219728
rect 76480 219320 77724 219321
rect 76480 218242 76989 219320
rect 77245 219319 77724 219320
rect 78756 216815 79191 219733
rect 98977 219728 101152 219750
rect 101273 219732 101691 219853
rect 123575 219839 123653 219896
rect 123878 219853 123971 220086
rect 145968 220086 145974 220103
rect 146038 220086 146046 220103
rect 145968 220077 146046 220086
rect 146076 220103 146154 220113
rect 146076 220086 146083 220103
rect 146147 220086 146154 220103
rect 146076 219916 146154 220086
rect 146578 220103 146666 220114
rect 146578 220086 146584 220103
rect 146659 220086 146666 220103
rect 146578 220081 146666 220086
rect 168468 220103 168546 220307
rect 168649 220183 170535 220203
rect 168649 220150 168657 220183
rect 168649 220148 168680 220150
rect 169445 220148 170535 220183
rect 168649 220141 170535 220148
rect 189967 220120 190046 220515
rect 208364 220483 211665 221021
rect 212245 220515 212675 221020
rect 208371 220365 208710 220483
rect 208371 220204 208568 220365
rect 192749 220203 193020 220204
rect 190171 220184 193020 220203
rect 190171 220150 190186 220184
rect 192127 220150 193020 220184
rect 190171 220141 193020 220150
rect 190171 220137 192166 220141
rect 208467 220136 208544 220204
rect 213649 220200 215511 220203
rect 208668 220183 218657 220200
rect 208668 220178 213657 220183
rect 213691 220178 218657 220183
rect 208668 220148 208679 220178
rect 218645 220148 218657 220178
rect 208668 220138 218657 220148
rect 208467 220133 208546 220136
rect 168468 220086 168474 220103
rect 168538 220086 168546 220103
rect 146075 219896 146154 219916
rect 123373 219771 123653 219839
rect 123373 219763 123652 219771
rect 122708 219762 123652 219763
rect 98977 219321 100949 219728
rect 101074 219725 101152 219728
rect 98977 218223 99481 219321
rect 99745 219319 100224 219321
rect 101256 216843 101691 219732
rect 121480 219728 123652 219762
rect 121480 219321 123449 219728
rect 123574 219725 123652 219728
rect 121480 219320 122724 219321
rect 121480 218165 121960 219320
rect 122245 219319 122724 219320
rect 123756 216846 124191 219853
rect 146075 219839 146153 219896
rect 146577 219853 146667 220081
rect 168468 220077 168546 220086
rect 168576 220103 168654 220113
rect 168576 220086 168583 220103
rect 168647 220086 168654 220103
rect 168576 219916 168654 220086
rect 169478 220103 169566 220114
rect 169478 220086 169484 220103
rect 169559 220086 169566 220103
rect 169478 220059 169566 220086
rect 189968 220103 190046 220120
rect 189968 220086 189974 220103
rect 190038 220086 190046 220103
rect 189968 220077 190046 220086
rect 190076 220103 190154 220113
rect 190076 220086 190083 220103
rect 190147 220086 190154 220103
rect 168575 219896 168654 219916
rect 169480 219896 169566 220059
rect 190076 219916 190154 220086
rect 192178 220103 192265 220114
rect 192178 220086 192184 220103
rect 192259 220086 192265 220103
rect 192178 220070 192265 220086
rect 208468 220103 208546 220133
rect 208468 220086 208474 220103
rect 208538 220086 208546 220103
rect 208468 220077 208546 220086
rect 208576 220103 208654 220113
rect 208576 220086 208583 220103
rect 208647 220086 208654 220103
rect 218678 220103 218766 220114
rect 218678 220099 218684 220103
rect 192178 220066 192266 220070
rect 190075 219896 190154 219916
rect 145873 219771 146153 219839
rect 145873 219763 146152 219771
rect 145208 219762 146152 219763
rect 143980 219728 146152 219762
rect 143980 219321 145949 219728
rect 146074 219725 146152 219728
rect 143980 219319 145224 219321
rect 143980 219318 144920 219319
rect 143980 218205 144484 219318
rect 33745 216420 34192 216632
rect 56240 216330 56696 216767
rect 78744 216612 79191 216815
rect 78744 216452 79192 216612
rect 101246 216602 101691 216843
rect 78744 216374 79179 216452
rect 101246 216218 101690 216602
rect 123738 216293 124200 216846
rect 146256 216624 146691 219853
rect 168575 219839 168653 219896
rect 168373 219771 168653 219839
rect 166480 219762 166985 219764
rect 168373 219763 168652 219771
rect 167708 219762 168652 219763
rect 166480 219728 168652 219762
rect 166480 219321 168449 219728
rect 168574 219725 168652 219728
rect 166480 219320 167724 219321
rect 166480 218244 166985 219320
rect 167245 219319 167724 219320
rect 146244 216458 146693 216624
rect 169435 216392 169912 219896
rect 190075 219869 190153 219896
rect 189429 219867 190153 219869
rect 188985 219734 190153 219867
rect 192177 219824 192266 220066
rect 208576 219916 208654 220086
rect 218677 220086 218684 220099
rect 218759 220086 218766 220103
rect 218677 219951 218766 220086
rect 208575 219896 208654 219916
rect 208575 219881 208653 219896
rect 208576 219865 208653 219881
rect 192177 219797 192267 219824
rect 188985 218027 189484 219734
rect 190075 219733 190153 219734
rect 192178 219606 192267 219797
rect 192177 219555 192267 219606
rect 192177 219132 192266 219555
rect 192177 219107 192267 219132
rect 192178 218904 192267 219107
rect 192104 216333 192426 218904
rect 208524 218238 208750 219865
rect 208524 217062 211612 218238
rect 208524 217056 208750 217062
rect 218625 217023 218871 219951
rect 215896 216737 218871 217023
rect 215896 215980 218864 216737
rect 10932 197349 11171 197645
rect 10968 197307 11045 197349
rect 10968 197103 11046 197307
rect 13010 197203 13515 197368
rect 33409 197355 33743 197714
rect 11149 197183 13515 197203
rect 11149 197150 11157 197183
rect 11191 197150 13515 197183
rect 11149 197141 13515 197150
rect 10968 197073 10974 197103
rect 11038 197073 11046 197103
rect 10968 197064 11046 197073
rect 11076 197103 11154 197113
rect 11076 197073 11083 197103
rect 11147 197073 11154 197103
rect 11076 196916 11154 197073
rect 11075 196896 11154 196916
rect 11193 197103 11281 197114
rect 11193 197073 11199 197103
rect 11274 197073 11281 197103
rect 11193 197061 11281 197073
rect 11075 196839 11153 196896
rect 10873 196771 11153 196839
rect 11193 196853 11271 197061
rect 11193 196802 11691 196853
rect 10873 196763 11152 196771
rect 10208 196762 11152 196763
rect 8981 196728 11152 196762
rect 11194 196733 11691 196802
rect 8981 196504 10949 196728
rect 11074 196725 11152 196728
rect 8980 196321 10949 196504
rect 8980 196319 10224 196321
rect 8980 195250 9482 196319
rect 8980 193650 9485 195250
rect 11256 194006 11691 196733
rect 13010 195755 13515 197141
rect 33468 197307 33545 197355
rect 33468 197103 33546 197307
rect 35510 197203 36015 197368
rect 55798 197325 56242 197641
rect 33649 197183 36015 197203
rect 33649 197150 33657 197183
rect 33691 197150 36015 197183
rect 33649 197141 36015 197150
rect 33468 197073 33474 197103
rect 33538 197073 33546 197103
rect 33468 197064 33546 197073
rect 33576 197103 33654 197113
rect 33576 197073 33583 197103
rect 33647 197073 33654 197103
rect 33576 196916 33654 197073
rect 33696 197103 33784 197114
rect 33696 197073 33702 197103
rect 33777 197073 33784 197103
rect 33696 197061 33784 197073
rect 33696 197059 33774 197061
rect 33696 197018 33771 197059
rect 33575 196896 33654 196916
rect 33575 196839 33653 196896
rect 33373 196771 33653 196839
rect 33693 196853 33771 197018
rect 33693 196802 34191 196853
rect 31479 196762 32255 196764
rect 33373 196763 33652 196771
rect 32708 196762 33652 196763
rect 31479 196728 33652 196762
rect 33694 196733 34191 196802
rect 31479 196321 33449 196728
rect 33574 196725 33652 196728
rect 31479 196319 32724 196321
rect 31479 195249 32255 196319
rect 11246 193261 11696 194006
rect 31480 193650 31985 195249
rect 33756 193747 34191 196733
rect 35510 195755 36015 197141
rect 55968 197103 56046 197325
rect 58010 197204 58515 197368
rect 78407 197351 78609 197561
rect 57750 197203 58515 197204
rect 56149 197183 58515 197203
rect 56149 197150 56157 197183
rect 56191 197150 58515 197183
rect 56149 197141 58515 197150
rect 55968 197073 55974 197103
rect 56038 197073 56046 197103
rect 55968 197064 56046 197073
rect 56076 197103 56154 197113
rect 56076 197073 56083 197103
rect 56147 197073 56154 197103
rect 56076 196916 56154 197073
rect 56075 196896 56154 196916
rect 56203 197103 56291 197114
rect 56203 197073 56209 197103
rect 56284 197073 56291 197103
rect 56203 197061 56291 197073
rect 56075 196839 56153 196896
rect 55873 196771 56153 196839
rect 56203 196853 56281 197061
rect 56203 196802 56691 196853
rect 55873 196763 56152 196771
rect 55208 196762 56152 196763
rect 53983 196755 54481 196761
rect 54745 196755 56152 196762
rect 53983 196728 56152 196755
rect 56204 196733 56691 196802
rect 53983 196327 55949 196728
rect 56074 196725 56152 196728
rect 56225 196626 56691 196733
rect 53983 195250 54481 196327
rect 54745 196321 55949 196327
rect 54745 196319 55224 196321
rect 33748 193431 34192 193747
rect 53980 193650 54485 195250
rect 56256 193767 56691 196626
rect 58010 195755 58515 197141
rect 78468 197307 78545 197351
rect 78468 197103 78546 197307
rect 80510 197203 81015 197368
rect 100788 197356 101240 197866
rect 78649 197183 81015 197203
rect 78649 197150 78657 197183
rect 78691 197150 81015 197183
rect 78649 197141 81015 197150
rect 78468 197073 78474 197103
rect 78538 197073 78546 197103
rect 78468 197064 78546 197073
rect 78576 197103 78654 197113
rect 78576 197073 78583 197103
rect 78647 197073 78654 197103
rect 78576 196916 78654 197073
rect 78575 196896 78654 196916
rect 78728 197103 78816 197114
rect 78728 197073 78734 197103
rect 78809 197073 78816 197103
rect 78728 197061 78816 197073
rect 78575 196839 78653 196896
rect 78373 196771 78653 196839
rect 78728 196853 78806 197061
rect 78728 196802 79191 196853
rect 76480 196761 76989 196764
rect 78373 196763 78652 196771
rect 77708 196762 78652 196763
rect 77245 196761 78652 196762
rect 76480 196728 78652 196761
rect 78729 196733 79191 196802
rect 76480 196321 78449 196728
rect 78574 196725 78652 196728
rect 76480 196320 77724 196321
rect 76480 195242 76989 196320
rect 77245 196319 77724 196320
rect 56240 193666 56696 193767
rect 56240 193650 56697 193666
rect 76480 193650 76985 195242
rect 78756 193815 79191 196733
rect 80510 195755 81015 197141
rect 100968 197307 101045 197356
rect 100968 197103 101046 197307
rect 103010 197203 103515 197368
rect 123259 197361 123733 197793
rect 101149 197183 103515 197203
rect 101149 197150 101157 197183
rect 101191 197150 103515 197183
rect 101149 197141 103515 197150
rect 100968 197073 100974 197103
rect 101038 197073 101046 197103
rect 100968 197064 101046 197073
rect 101076 197103 101154 197113
rect 101076 197073 101083 197103
rect 101147 197073 101154 197103
rect 101076 196916 101154 197073
rect 101278 197103 101366 197114
rect 101278 197073 101284 197103
rect 101359 197073 101366 197103
rect 101278 197061 101366 197073
rect 101278 197031 101356 197061
rect 101075 196896 101154 196916
rect 101075 196839 101153 196896
rect 101277 196853 101357 197031
rect 100873 196771 101153 196839
rect 100873 196763 101152 196771
rect 100208 196762 101152 196763
rect 99745 196760 101152 196762
rect 99230 196750 101152 196760
rect 98977 196728 101152 196750
rect 101273 196732 101691 196853
rect 98977 196321 100949 196728
rect 101074 196725 101152 196728
rect 98977 195250 99481 196321
rect 99745 196319 100224 196321
rect 98977 195223 99485 195250
rect 78744 193650 79191 193815
rect 98980 193650 99485 195223
rect 101256 193843 101691 196732
rect 103010 195755 103515 197141
rect 123468 197307 123545 197361
rect 123468 197103 123546 197307
rect 125510 197203 126015 197368
rect 145793 197353 146245 197801
rect 123649 197183 126015 197203
rect 123649 197150 123657 197183
rect 123649 197149 123691 197150
rect 123860 197149 126015 197183
rect 123649 197141 126015 197149
rect 125242 197140 126015 197141
rect 123468 197073 123474 197103
rect 123538 197073 123546 197103
rect 123468 197064 123546 197073
rect 123576 197103 123654 197113
rect 123576 197073 123583 197103
rect 123647 197073 123654 197103
rect 123576 196916 123654 197073
rect 123575 196896 123654 196916
rect 123878 197103 123966 197114
rect 123878 197073 123884 197103
rect 123959 197098 123966 197103
rect 123959 197073 123971 197098
rect 123575 196839 123653 196896
rect 123878 196853 123971 197073
rect 123373 196771 123653 196839
rect 123373 196763 123652 196771
rect 122708 196762 123652 196763
rect 121480 196728 123652 196762
rect 121480 196321 123449 196728
rect 123574 196725 123652 196728
rect 121480 196320 122724 196321
rect 101246 193840 101691 193843
rect 121480 195250 121960 196320
rect 122245 196319 122724 196320
rect 56253 193350 56697 193650
rect 78748 193455 79189 193650
rect 101246 193330 101698 193840
rect 121480 193650 121985 195250
rect 123756 193846 124191 196853
rect 125510 195755 126015 197140
rect 145968 197307 146045 197353
rect 145968 197103 146046 197307
rect 148010 197203 148515 197368
rect 168223 197357 168724 197817
rect 146149 197183 148515 197203
rect 146149 197150 146157 197183
rect 146149 197148 146178 197150
rect 146552 197148 148515 197183
rect 146149 197141 148515 197148
rect 145968 197073 145974 197103
rect 146038 197073 146046 197103
rect 145968 197064 146046 197073
rect 146076 197103 146154 197113
rect 146076 197073 146083 197103
rect 146147 197073 146154 197103
rect 146578 197103 146666 197114
rect 146578 197081 146584 197103
rect 146076 196916 146154 197073
rect 146075 196896 146154 196916
rect 146577 197073 146584 197081
rect 146659 197081 146666 197103
rect 146659 197073 146667 197081
rect 146075 196839 146153 196896
rect 146577 196853 146667 197073
rect 145873 196771 146153 196839
rect 145873 196763 146152 196771
rect 145208 196762 146152 196763
rect 143980 196728 146152 196762
rect 143980 196321 145949 196728
rect 146074 196725 146152 196728
rect 143980 196319 145224 196321
rect 143980 196318 144920 196319
rect 143980 195250 144484 196318
rect 123738 193773 124200 193846
rect 123738 193650 124219 193773
rect 143980 193650 144485 195250
rect 146256 193693 146691 196853
rect 148010 195755 148515 197141
rect 168468 197307 168545 197357
rect 168468 197103 168546 197307
rect 170510 197203 171015 197368
rect 189837 197367 190147 197928
rect 208436 197726 211959 198016
rect 208371 197515 211959 197726
rect 168649 197183 171015 197203
rect 168649 197150 168657 197183
rect 168649 197148 168680 197150
rect 169445 197148 171015 197183
rect 168649 197141 171015 197148
rect 168468 197073 168474 197103
rect 168538 197073 168546 197103
rect 168468 197064 168546 197073
rect 168576 197103 168654 197113
rect 168576 197073 168583 197103
rect 168647 197073 168654 197103
rect 168576 196916 168654 197073
rect 169478 197103 169566 197114
rect 169478 197073 169484 197103
rect 169559 197073 169566 197103
rect 169478 197059 169566 197073
rect 168575 196896 168654 196916
rect 169480 196896 169566 197059
rect 168575 196839 168653 196896
rect 168373 196771 168653 196839
rect 166480 196762 166985 196764
rect 168373 196763 168652 196771
rect 167708 196762 168652 196763
rect 166480 196728 168652 196762
rect 166480 196321 168449 196728
rect 168574 196725 168652 196728
rect 166480 196320 167724 196321
rect 146256 193650 146709 193693
rect 166480 193650 166985 196320
rect 167245 196319 167724 196320
rect 169435 193791 169912 196896
rect 170510 195755 171015 197141
rect 189967 197120 190046 197367
rect 193010 197204 193515 197368
rect 208371 197367 208827 197515
rect 208371 197365 208710 197367
rect 208371 197204 208568 197365
rect 192749 197203 193515 197204
rect 190171 197184 193515 197203
rect 190171 197150 190186 197184
rect 192127 197150 193515 197184
rect 190171 197141 193515 197150
rect 190171 197137 192166 197141
rect 189968 197103 190046 197120
rect 189968 197073 189974 197103
rect 190038 197073 190046 197103
rect 189968 197064 190046 197073
rect 190076 197103 190154 197113
rect 190076 197073 190083 197103
rect 190147 197073 190154 197103
rect 190076 196916 190154 197073
rect 192178 197103 192266 197114
rect 192178 197073 192184 197103
rect 192259 197073 192266 197103
rect 192178 197066 192266 197073
rect 190075 196896 190154 196916
rect 190075 196869 190153 196896
rect 189429 196867 190153 196869
rect 188985 196734 190153 196867
rect 192177 196824 192266 197066
rect 192177 196797 192267 196824
rect 188985 195250 189484 196734
rect 190075 196733 190153 196734
rect 192178 196606 192267 196797
rect 192177 196555 192267 196606
rect 192177 196132 192266 196555
rect 192177 196107 192267 196132
rect 192178 195904 192267 196107
rect 123745 193341 124219 193650
rect 146257 193245 146709 193650
rect 169418 193331 169919 193791
rect 188980 193650 189485 195250
rect 192104 194023 192426 195904
rect 193010 195755 193515 197141
rect 208467 197136 208544 197204
rect 215510 197203 216015 197368
rect 213649 197200 216015 197203
rect 208668 197183 218657 197200
rect 208668 197178 213657 197183
rect 213691 197178 218657 197183
rect 208668 197148 208679 197178
rect 218645 197148 218657 197178
rect 208668 197138 218657 197148
rect 208467 197133 208546 197136
rect 208468 197103 208546 197133
rect 208468 197073 208474 197103
rect 208538 197073 208546 197103
rect 208468 197064 208546 197073
rect 208576 197103 208654 197113
rect 208576 197073 208583 197103
rect 208647 197073 208654 197103
rect 208576 196916 208654 197073
rect 208575 196896 208654 196916
rect 208575 196881 208653 196896
rect 208576 196865 208653 196881
rect 208524 195238 208750 196865
rect 215510 195755 216015 197138
rect 218678 197103 218766 197114
rect 218678 197099 218684 197103
rect 218677 197073 218684 197099
rect 218759 197073 218766 197103
rect 218677 196951 218766 197073
rect 211480 195238 211985 195250
rect 208524 194062 211985 195238
rect 208524 194056 208750 194062
rect 192104 193650 192427 194023
rect 211480 193650 211985 194062
rect 218625 194023 218871 196951
rect 215896 193737 218871 194023
rect 215896 193650 218864 193737
rect 192109 193266 192427 193650
rect 55659 174826 56107 174866
rect 168286 174827 168734 174832
rect 10868 174366 11250 174770
rect 10968 174307 11045 174366
rect 10968 174103 11046 174307
rect 13010 174203 13515 174368
rect 33291 174354 33739 174814
rect 55659 174406 56212 174826
rect 11149 174183 13515 174203
rect 11149 174150 11157 174183
rect 11191 174150 13515 174183
rect 11149 174141 13515 174150
rect 10968 174064 10974 174103
rect 11038 174064 11046 174103
rect 10968 174055 11046 174064
rect 11076 174103 11154 174113
rect 11076 174064 11083 174103
rect 11147 174064 11154 174103
rect 11076 173916 11154 174064
rect 11075 173896 11154 173916
rect 11193 174103 11281 174114
rect 11193 174064 11199 174103
rect 11274 174064 11281 174103
rect 11193 174052 11281 174064
rect 11075 173839 11153 173896
rect 10873 173771 11153 173839
rect 11193 173853 11271 174052
rect 11193 173802 11691 173853
rect 10873 173763 11152 173771
rect 10208 173762 11152 173763
rect 8981 173728 11152 173762
rect 11194 173733 11691 173802
rect 8981 173504 10949 173728
rect 11074 173725 11152 173728
rect 8980 173321 10949 173504
rect 8980 173319 10224 173321
rect 8980 172250 9482 173319
rect 8980 170650 9485 172250
rect 11256 170790 11691 173733
rect 13010 172755 13515 174141
rect 33468 174307 33545 174354
rect 33468 174103 33546 174307
rect 35510 174203 36015 174368
rect 55764 174366 56212 174406
rect 33649 174183 36015 174203
rect 33649 174150 33657 174183
rect 33691 174150 36015 174183
rect 33649 174141 36015 174150
rect 33468 174064 33474 174103
rect 33538 174064 33546 174103
rect 33468 174055 33546 174064
rect 33576 174103 33654 174113
rect 33576 174064 33583 174103
rect 33647 174064 33654 174103
rect 33576 173916 33654 174064
rect 33696 174103 33784 174114
rect 33696 174064 33702 174103
rect 33777 174064 33784 174103
rect 33696 174052 33784 174064
rect 33696 174018 33771 174052
rect 33575 173896 33654 173916
rect 33575 173839 33653 173896
rect 33373 173771 33653 173839
rect 33693 173853 33771 174018
rect 33693 173802 34191 173853
rect 31479 173762 32255 173764
rect 33373 173763 33652 173771
rect 32708 173762 33652 173763
rect 31479 173728 33652 173762
rect 33694 173733 34191 173802
rect 31479 173321 33449 173728
rect 33574 173725 33652 173728
rect 31479 173319 32724 173321
rect 31479 172249 32255 173319
rect 11245 170330 11693 170790
rect 31480 170650 31985 172249
rect 33756 170780 34191 173733
rect 35510 172755 36015 174141
rect 55968 174307 56045 174366
rect 55968 174103 56046 174307
rect 58010 174204 58515 174368
rect 78301 174364 78749 174824
rect 57750 174203 58515 174204
rect 56149 174183 58515 174203
rect 56149 174150 56157 174183
rect 56191 174150 58515 174183
rect 56149 174141 58515 174150
rect 55968 174064 55974 174103
rect 56038 174064 56046 174103
rect 55968 174055 56046 174064
rect 56076 174103 56154 174113
rect 56076 174064 56083 174103
rect 56147 174064 56154 174103
rect 56076 173916 56154 174064
rect 56075 173896 56154 173916
rect 56203 174103 56291 174114
rect 56203 174064 56209 174103
rect 56284 174064 56291 174103
rect 56203 174052 56291 174064
rect 56075 173839 56153 173896
rect 55873 173771 56153 173839
rect 56203 173853 56281 174052
rect 56203 173802 56691 173853
rect 55873 173763 56152 173771
rect 55208 173762 56152 173763
rect 53983 173755 54481 173761
rect 54745 173755 56152 173762
rect 53983 173728 56152 173755
rect 56204 173733 56691 173802
rect 53983 173327 55949 173728
rect 56074 173725 56152 173728
rect 56225 173626 56691 173733
rect 53983 172250 54481 173327
rect 54745 173321 55949 173327
rect 54745 173319 55224 173321
rect 33745 170320 34193 170780
rect 53980 170650 54485 172250
rect 56256 170767 56691 173626
rect 58010 172755 58515 174141
rect 78468 174307 78545 174364
rect 78468 174103 78546 174307
rect 80510 174203 81015 174368
rect 100761 174360 101209 174820
rect 78649 174183 81015 174203
rect 78649 174150 78657 174183
rect 78691 174150 81015 174183
rect 78649 174141 81015 174150
rect 78468 174064 78474 174103
rect 78538 174064 78546 174103
rect 78468 174055 78546 174064
rect 78576 174103 78654 174113
rect 78576 174064 78583 174103
rect 78647 174064 78654 174103
rect 78576 173916 78654 174064
rect 78575 173896 78654 173916
rect 78728 174103 78816 174114
rect 78728 174064 78734 174103
rect 78809 174064 78816 174103
rect 78728 174052 78816 174064
rect 78575 173839 78653 173896
rect 78373 173771 78653 173839
rect 78728 173853 78806 174052
rect 78728 173802 79191 173853
rect 76480 173761 76989 173764
rect 78373 173763 78652 173771
rect 77708 173762 78652 173763
rect 77245 173761 78652 173762
rect 76480 173728 78652 173761
rect 78729 173733 79191 173802
rect 76480 173321 78449 173728
rect 78574 173725 78652 173728
rect 76480 173320 77724 173321
rect 76480 172242 76989 173320
rect 77245 173319 77724 173320
rect 56240 170661 56696 170767
rect 56227 170650 56696 170661
rect 76480 170650 76985 172242
rect 78756 170895 79191 173733
rect 80510 172755 81015 174141
rect 100968 174307 101045 174360
rect 100968 174103 101046 174307
rect 103010 174203 103515 174368
rect 123281 174363 123729 174823
rect 101149 174183 103515 174203
rect 101149 174150 101157 174183
rect 101191 174150 103515 174183
rect 101149 174141 103515 174150
rect 100968 174064 100974 174103
rect 101038 174064 101046 174103
rect 100968 174055 101046 174064
rect 101076 174103 101154 174113
rect 101076 174064 101083 174103
rect 101147 174064 101154 174103
rect 101076 173916 101154 174064
rect 101278 174103 101366 174114
rect 101278 174064 101284 174103
rect 101359 174064 101366 174103
rect 101278 174052 101366 174064
rect 101278 174031 101356 174052
rect 101075 173896 101154 173916
rect 101075 173839 101153 173896
rect 101277 173853 101357 174031
rect 100873 173771 101153 173839
rect 100873 173763 101152 173771
rect 100208 173762 101152 173763
rect 99745 173760 101152 173762
rect 99230 173750 101152 173760
rect 98977 173728 101152 173750
rect 101273 173732 101691 173853
rect 98977 173321 100949 173728
rect 101074 173725 101152 173728
rect 98977 172250 99481 173321
rect 99745 173319 100224 173321
rect 98977 172223 99485 172250
rect 78740 170650 79191 170895
rect 98980 170650 99485 172223
rect 101256 170843 101691 173732
rect 103010 172755 103515 174141
rect 123468 174307 123545 174363
rect 123468 174103 123546 174307
rect 125510 174203 126015 174368
rect 145762 174360 146210 174820
rect 168280 174372 168734 174827
rect 123649 174183 126015 174203
rect 123649 174150 123657 174183
rect 123649 174149 123691 174150
rect 123860 174149 126015 174183
rect 123649 174141 126015 174149
rect 125242 174140 126015 174141
rect 123468 174064 123474 174103
rect 123538 174064 123546 174103
rect 123468 174055 123546 174064
rect 123576 174103 123654 174113
rect 123576 174064 123583 174103
rect 123647 174064 123654 174103
rect 123576 173916 123654 174064
rect 123575 173896 123654 173916
rect 123878 174103 123966 174114
rect 123878 174064 123884 174103
rect 123959 174098 123966 174103
rect 123959 174064 123971 174098
rect 123575 173839 123653 173896
rect 123878 173853 123971 174064
rect 123373 173771 123653 173839
rect 123373 173763 123652 173771
rect 122708 173762 123652 173763
rect 121480 173728 123652 173762
rect 121480 173321 123449 173728
rect 123574 173725 123652 173728
rect 121480 173320 122724 173321
rect 101246 170842 101691 170843
rect 101232 170650 101691 170842
rect 121480 172250 121960 173320
rect 122245 173319 122724 173320
rect 121480 170650 121985 172250
rect 123756 170931 124191 173853
rect 125510 172755 126015 174140
rect 145968 174307 146045 174360
rect 145968 174103 146046 174307
rect 148010 174203 148515 174368
rect 168280 174367 168728 174372
rect 189764 174368 190212 174828
rect 208580 174825 211596 175022
rect 208357 174522 211596 174825
rect 146149 174183 148515 174203
rect 146149 174150 146157 174183
rect 146149 174148 146178 174150
rect 146552 174148 148515 174183
rect 146149 174141 148515 174148
rect 145968 174064 145974 174103
rect 146038 174064 146046 174103
rect 145968 174055 146046 174064
rect 146076 174103 146154 174113
rect 146076 174064 146083 174103
rect 146147 174064 146154 174103
rect 146578 174103 146666 174114
rect 146578 174081 146584 174103
rect 146076 173916 146154 174064
rect 146075 173896 146154 173916
rect 146577 174064 146584 174081
rect 146659 174081 146666 174103
rect 146659 174064 146667 174081
rect 146075 173839 146153 173896
rect 146577 173853 146667 174064
rect 145873 173771 146153 173839
rect 145873 173763 146152 173771
rect 145208 173762 146152 173763
rect 143980 173728 146152 173762
rect 143980 173321 145949 173728
rect 146074 173725 146152 173728
rect 143980 173319 145224 173321
rect 143980 173318 144920 173319
rect 143980 172250 144484 173318
rect 123745 170846 124193 170931
rect 123738 170650 124200 170846
rect 143980 170650 144485 172250
rect 146256 170837 146691 173853
rect 148010 172755 148515 174141
rect 168468 174307 168545 174367
rect 168468 174103 168546 174307
rect 170510 174203 171015 174368
rect 168649 174183 171015 174203
rect 168649 174150 168657 174183
rect 168649 174148 168680 174150
rect 169445 174148 171015 174183
rect 168649 174141 171015 174148
rect 168468 174064 168474 174103
rect 168538 174064 168546 174103
rect 168468 174055 168546 174064
rect 168576 174103 168654 174113
rect 168576 174064 168583 174103
rect 168647 174064 168654 174103
rect 168576 173916 168654 174064
rect 169478 174103 169566 174114
rect 169478 174064 169484 174103
rect 169559 174064 169566 174103
rect 169478 174052 169566 174064
rect 168575 173896 168654 173916
rect 169480 173896 169566 174052
rect 168575 173839 168653 173896
rect 168373 173771 168653 173839
rect 166480 173762 166985 173764
rect 168373 173763 168652 173771
rect 167708 173762 168652 173763
rect 166480 173728 168652 173762
rect 166480 173321 168449 173728
rect 168574 173725 168652 173728
rect 166480 173320 167724 173321
rect 146232 170650 146691 170837
rect 166480 170650 166985 173320
rect 167245 173319 167724 173320
rect 169435 170650 169912 173896
rect 170510 172755 171015 174141
rect 189967 174120 190046 174368
rect 193010 174204 193515 174368
rect 208357 174365 208805 174522
rect 208371 174204 208568 174365
rect 192749 174203 193515 174204
rect 190171 174184 193515 174203
rect 190171 174150 190186 174184
rect 192127 174150 193515 174184
rect 190171 174141 193515 174150
rect 190171 174137 192166 174141
rect 189968 174103 190046 174120
rect 189968 174064 189974 174103
rect 190038 174064 190046 174103
rect 189968 174055 190046 174064
rect 190076 174103 190154 174113
rect 190076 174064 190083 174103
rect 190147 174064 190154 174103
rect 192178 174103 192266 174114
rect 192178 174066 192184 174103
rect 190076 173916 190154 174064
rect 190075 173896 190154 173916
rect 192177 174064 192184 174066
rect 192259 174064 192266 174103
rect 190075 173869 190153 173896
rect 189429 173867 190153 173869
rect 188985 173734 190153 173867
rect 192177 173824 192266 174064
rect 192177 173797 192267 173824
rect 188985 172250 189484 173734
rect 190075 173733 190153 173734
rect 192178 173606 192267 173797
rect 192177 173555 192267 173606
rect 192177 173132 192266 173555
rect 192177 173107 192267 173132
rect 192178 172904 192267 173107
rect 188980 170650 189485 172250
rect 192104 170830 192426 172904
rect 193010 172755 193515 174141
rect 208467 174136 208544 174204
rect 215510 174203 216015 174368
rect 213649 174200 216015 174203
rect 208668 174183 218657 174200
rect 208668 174178 213657 174183
rect 213691 174178 218657 174183
rect 208668 174148 208679 174178
rect 218645 174148 218657 174178
rect 208668 174138 218657 174148
rect 208467 174133 208546 174136
rect 208468 174103 208546 174133
rect 208468 174064 208474 174103
rect 208538 174064 208546 174103
rect 208468 174055 208546 174064
rect 208576 174103 208654 174113
rect 208576 174064 208583 174103
rect 208647 174064 208654 174103
rect 208576 173916 208654 174064
rect 208575 173896 208654 173916
rect 208575 173881 208653 173896
rect 208576 173865 208653 173881
rect 208524 172238 208750 173865
rect 215510 172755 216015 174138
rect 218678 174103 218766 174114
rect 218678 174099 218684 174103
rect 218677 174064 218684 174099
rect 218759 174064 218766 174103
rect 218677 173951 218766 174064
rect 211480 172238 211985 172250
rect 208524 171062 211985 172238
rect 208524 171056 208750 171062
rect 56227 170201 56675 170650
rect 78740 170435 79188 170650
rect 101232 170382 101680 170650
rect 123745 170471 124193 170650
rect 146232 170377 146680 170650
rect 169439 170289 169887 170650
rect 192069 170370 192517 170830
rect 211480 170650 211985 171062
rect 215510 171023 216010 171025
rect 218625 171023 218871 173951
rect 215510 170737 218871 171023
rect 215510 170650 218864 170737
rect 215510 169975 216010 170650
rect 208262 152372 209925 152400
rect 78258 152246 78725 152252
rect 10796 151364 11257 152111
rect 10968 151307 11045 151364
rect 10968 151103 11046 151307
rect 13010 151203 13515 151368
rect 33312 151357 33719 151912
rect 55906 151368 56246 151572
rect 78258 151371 78726 152246
rect 100900 151982 101231 152005
rect 11149 151183 13515 151203
rect 11149 151150 11157 151183
rect 11191 151150 13515 151183
rect 11149 151141 13515 151150
rect 10968 151044 10974 151103
rect 11038 151044 11046 151103
rect 10968 151035 11046 151044
rect 11076 151103 11154 151113
rect 11076 151044 11083 151103
rect 11147 151044 11154 151103
rect 11076 150916 11154 151044
rect 11075 150896 11154 150916
rect 11193 151103 11281 151114
rect 11193 151044 11199 151103
rect 11274 151044 11281 151103
rect 11193 151032 11281 151044
rect 11075 150839 11153 150896
rect 10873 150771 11153 150839
rect 11193 150853 11271 151032
rect 11193 150802 11691 150853
rect 10873 150763 11152 150771
rect 10208 150762 11152 150763
rect 8981 150728 11152 150762
rect 11194 150733 11691 150802
rect 8981 150504 10949 150728
rect 11074 150725 11152 150728
rect 8980 150321 10949 150504
rect 8980 150319 10224 150321
rect 8980 149250 9482 150319
rect 8980 147650 9485 149250
rect 11256 147919 11691 150733
rect 13010 149755 13515 151141
rect 33468 151307 33545 151357
rect 33468 151103 33546 151307
rect 35510 151203 36015 151368
rect 33649 151183 36015 151203
rect 33649 151150 33657 151183
rect 33691 151150 36015 151183
rect 33649 151141 36015 151150
rect 33468 151044 33474 151103
rect 33538 151044 33546 151103
rect 33468 151035 33546 151044
rect 33576 151103 33654 151113
rect 33576 151044 33583 151103
rect 33647 151044 33654 151103
rect 33576 150916 33654 151044
rect 33696 151103 33784 151114
rect 33696 151044 33702 151103
rect 33777 151044 33784 151103
rect 33696 151032 33784 151044
rect 33696 151018 33771 151032
rect 33575 150896 33654 150916
rect 33575 150839 33653 150896
rect 33373 150771 33653 150839
rect 33693 150853 33771 151018
rect 33693 150802 34191 150853
rect 31479 150762 32255 150764
rect 33373 150763 33652 150771
rect 32708 150762 33652 150763
rect 31479 150728 33652 150762
rect 33694 150733 34191 150802
rect 31479 150321 33449 150728
rect 33574 150725 33652 150728
rect 31479 150319 32724 150321
rect 31479 149249 32255 150319
rect 11246 147172 11707 147919
rect 31480 147650 31985 149249
rect 33756 147940 34191 150733
rect 35510 149755 36015 151141
rect 55968 151307 56045 151368
rect 55968 151103 56046 151307
rect 58010 151204 58515 151368
rect 78259 151365 78726 151371
rect 100894 151373 101231 151982
rect 57750 151203 58515 151204
rect 56149 151183 58515 151203
rect 56149 151150 56157 151183
rect 56191 151150 58515 151183
rect 56149 151141 58515 151150
rect 55968 151044 55974 151103
rect 56038 151044 56046 151103
rect 55968 151035 56046 151044
rect 56076 151103 56154 151113
rect 56076 151044 56083 151103
rect 56147 151044 56154 151103
rect 56076 150916 56154 151044
rect 56075 150896 56154 150916
rect 56203 151103 56291 151114
rect 56203 151044 56209 151103
rect 56284 151044 56291 151103
rect 56203 151032 56291 151044
rect 56075 150839 56153 150896
rect 55873 150771 56153 150839
rect 56203 150853 56281 151032
rect 56203 150802 56691 150853
rect 55873 150763 56152 150771
rect 55208 150762 56152 150763
rect 53983 150755 54481 150761
rect 54745 150755 56152 150762
rect 53983 150728 56152 150755
rect 56204 150733 56691 150802
rect 53983 150327 55949 150728
rect 56074 150725 56152 150728
rect 56225 150626 56691 150733
rect 53983 149250 54481 150327
rect 54745 150321 55949 150327
rect 54745 150319 55224 150321
rect 33738 147215 34193 147940
rect 53980 147650 54485 149250
rect 56256 148022 56691 150626
rect 58010 149755 58515 151141
rect 78468 151307 78545 151365
rect 78468 151103 78546 151307
rect 80510 151203 81015 151368
rect 100894 151350 101225 151373
rect 78649 151183 81015 151203
rect 78649 151150 78657 151183
rect 78691 151150 81015 151183
rect 78649 151141 81015 151150
rect 78468 151044 78474 151103
rect 78538 151044 78546 151103
rect 78468 151035 78546 151044
rect 78576 151103 78654 151113
rect 78576 151044 78583 151103
rect 78647 151044 78654 151103
rect 78576 150916 78654 151044
rect 78575 150896 78654 150916
rect 78728 151103 78816 151114
rect 78728 151044 78734 151103
rect 78809 151044 78816 151103
rect 78728 151032 78816 151044
rect 78575 150839 78653 150896
rect 78373 150771 78653 150839
rect 78728 150853 78806 151032
rect 78728 150802 79191 150853
rect 76480 150761 76989 150764
rect 78373 150763 78652 150771
rect 77708 150762 78652 150763
rect 77245 150761 78652 150762
rect 76480 150728 78652 150761
rect 78729 150733 79191 150802
rect 76480 150321 78449 150728
rect 78574 150725 78652 150728
rect 76480 150320 77724 150321
rect 76480 149242 76989 150320
rect 77245 150319 77724 150320
rect 56229 147767 56693 148022
rect 56229 147650 56696 147767
rect 76480 147650 76985 149242
rect 78756 148061 79191 150733
rect 80510 149755 81015 151141
rect 100968 151307 101045 151350
rect 100968 151103 101046 151307
rect 103010 151203 103515 151368
rect 123165 151352 123627 152033
rect 208262 152018 209926 152372
rect 145856 151368 146232 151719
rect 101149 151183 103515 151203
rect 101149 151150 101157 151183
rect 101191 151150 103515 151183
rect 101149 151141 103515 151150
rect 100968 151044 100974 151103
rect 101038 151044 101046 151103
rect 100968 151035 101046 151044
rect 101076 151103 101154 151113
rect 101076 151044 101083 151103
rect 101147 151044 101154 151103
rect 101076 150916 101154 151044
rect 101278 151103 101366 151114
rect 101278 151044 101284 151103
rect 101359 151044 101366 151103
rect 101278 151032 101366 151044
rect 101278 151031 101364 151032
rect 101075 150896 101154 150916
rect 101277 151015 101364 151031
rect 101075 150839 101153 150896
rect 101277 150853 101357 151015
rect 100873 150771 101153 150839
rect 100873 150763 101152 150771
rect 100208 150762 101152 150763
rect 99745 150760 101152 150762
rect 99230 150750 101152 150760
rect 98977 150728 101152 150750
rect 101273 150732 101691 150853
rect 98977 150321 100949 150728
rect 101074 150725 101152 150728
rect 98977 149250 99481 150321
rect 99745 150319 100224 150321
rect 98977 149223 99485 149250
rect 78746 147815 79213 148061
rect 78744 147650 79213 147815
rect 98980 147650 99485 149223
rect 101256 147966 101691 150732
rect 103010 149755 103515 151141
rect 123468 151307 123545 151352
rect 123468 151103 123546 151307
rect 125510 151203 126015 151368
rect 123649 151183 126015 151203
rect 123649 151150 123657 151183
rect 123649 151149 123691 151150
rect 123860 151149 126015 151183
rect 123649 151141 126015 151149
rect 125242 151140 126015 151141
rect 123468 151044 123474 151103
rect 123538 151044 123546 151103
rect 123468 151035 123546 151044
rect 123576 151103 123654 151113
rect 123576 151044 123583 151103
rect 123647 151044 123654 151103
rect 123576 150916 123654 151044
rect 123575 150896 123654 150916
rect 123878 151103 123966 151114
rect 123878 151044 123884 151103
rect 123959 151098 123966 151103
rect 123959 151044 123971 151098
rect 123575 150839 123653 150896
rect 123878 150853 123971 151044
rect 123373 150771 123653 150839
rect 123373 150763 123652 150771
rect 122708 150762 123652 150763
rect 121480 150728 123652 150762
rect 121480 150321 123449 150728
rect 123574 150725 123652 150728
rect 121480 150320 122724 150321
rect 121480 149250 121960 150320
rect 122245 150319 122724 150320
rect 56229 147223 56693 147650
rect 78746 147180 79213 147650
rect 101223 146997 101724 147966
rect 121480 147650 121985 149250
rect 123756 147946 124191 150853
rect 125510 149755 126015 151140
rect 145968 151307 146045 151368
rect 145968 151103 146046 151307
rect 148010 151203 148515 151368
rect 168311 151362 168743 151639
rect 146149 151183 148515 151203
rect 146149 151150 146157 151183
rect 146149 151148 146178 151150
rect 146552 151148 148515 151183
rect 146149 151141 148515 151148
rect 145968 151044 145974 151103
rect 146038 151044 146046 151103
rect 145968 151035 146046 151044
rect 146076 151103 146154 151113
rect 146076 151044 146083 151103
rect 146147 151044 146154 151103
rect 146578 151103 146666 151114
rect 146578 151081 146584 151103
rect 146076 150916 146154 151044
rect 146075 150896 146154 150916
rect 146577 151044 146584 151081
rect 146659 151081 146666 151103
rect 146659 151044 146667 151081
rect 146075 150839 146153 150896
rect 146577 150853 146667 151044
rect 145873 150771 146153 150839
rect 145873 150763 146152 150771
rect 145208 150762 146152 150763
rect 143980 150728 146152 150762
rect 143980 150321 145949 150728
rect 146074 150725 146152 150728
rect 143980 150319 145224 150321
rect 143980 150318 144920 150319
rect 143980 149250 144484 150318
rect 123756 147846 124220 147946
rect 123738 147650 124220 147846
rect 143980 147650 144485 149250
rect 146256 148078 146691 150853
rect 148010 149755 148515 151141
rect 168468 151307 168545 151362
rect 168468 151103 168546 151307
rect 170510 151203 171015 151368
rect 189809 151362 190194 151874
rect 208262 151527 211578 152018
rect 208262 151379 209926 151527
rect 168649 151183 171015 151203
rect 168649 151150 168657 151183
rect 168649 151148 168680 151150
rect 169445 151148 171015 151183
rect 168649 151141 171015 151148
rect 168468 151044 168474 151103
rect 168538 151044 168546 151103
rect 168468 151035 168546 151044
rect 168576 151103 168654 151113
rect 168576 151044 168583 151103
rect 168647 151044 168654 151103
rect 168576 150916 168654 151044
rect 169478 151103 169566 151114
rect 169478 151044 169484 151103
rect 169559 151044 169566 151103
rect 169478 151032 169566 151044
rect 168575 150896 168654 150916
rect 169480 150896 169566 151032
rect 168575 150839 168653 150896
rect 168373 150771 168653 150839
rect 166480 150762 166985 150764
rect 168373 150763 168652 150771
rect 167708 150762 168652 150763
rect 166480 150728 168652 150762
rect 166480 150321 168449 150728
rect 168574 150725 168652 150728
rect 166480 150320 167724 150321
rect 123758 147295 124220 147650
rect 146204 146975 146691 148078
rect 166480 147650 166985 150320
rect 167245 150319 167724 150320
rect 169435 147783 169912 150896
rect 170510 149755 171015 151141
rect 189967 151120 190046 151362
rect 193010 151204 193515 151368
rect 208263 151351 209926 151379
rect 208371 151204 208568 151351
rect 192749 151203 193515 151204
rect 190171 151184 193515 151203
rect 190171 151150 190186 151184
rect 192127 151150 193515 151184
rect 190171 151141 193515 151150
rect 190171 151137 192166 151141
rect 189968 151103 190046 151120
rect 189968 151044 189974 151103
rect 190038 151044 190046 151103
rect 189968 151035 190046 151044
rect 190076 151103 190154 151113
rect 190076 151044 190083 151103
rect 190147 151044 190154 151103
rect 192178 151103 192266 151114
rect 192178 151066 192184 151103
rect 190076 150916 190154 151044
rect 190075 150896 190154 150916
rect 192177 151044 192184 151066
rect 192259 151044 192266 151103
rect 190075 150869 190153 150896
rect 189429 150867 190153 150869
rect 188985 150734 190153 150867
rect 192177 150824 192266 151044
rect 192177 150797 192267 150824
rect 188985 149250 189484 150734
rect 190075 150733 190153 150734
rect 192178 150606 192267 150797
rect 192177 150555 192267 150606
rect 192177 150132 192266 150555
rect 192177 150107 192267 150132
rect 192178 149904 192267 150107
rect 169435 147650 169929 147783
rect 188980 147650 189485 149250
rect 192104 148155 192426 149904
rect 193010 149755 193515 151141
rect 208467 151136 208544 151204
rect 215510 151203 216015 151368
rect 213649 151200 216015 151203
rect 208668 151183 218657 151200
rect 208668 151178 213657 151183
rect 213691 151178 218657 151183
rect 208668 151148 208679 151178
rect 218645 151148 218657 151178
rect 208668 151138 218657 151148
rect 208467 151133 208546 151136
rect 208468 151103 208546 151133
rect 208468 151044 208474 151103
rect 208538 151044 208546 151103
rect 208468 151035 208546 151044
rect 208576 151103 208654 151113
rect 208576 151044 208583 151103
rect 208647 151044 208654 151103
rect 208576 150916 208654 151044
rect 208575 150896 208654 150916
rect 208575 150881 208653 150896
rect 208576 150865 208653 150881
rect 208524 149238 208750 150865
rect 215510 149755 216015 151138
rect 218678 151103 218766 151114
rect 218678 151099 218684 151103
rect 218677 151044 218684 151099
rect 218759 151044 218766 151103
rect 218677 150951 218766 151044
rect 211480 149238 211985 149250
rect 169438 147399 169929 147650
rect 192095 147258 192431 148155
rect 208524 148062 211985 149238
rect 208524 148056 208750 148062
rect 211480 147650 211985 148062
rect 215198 148023 216861 148024
rect 218625 148023 218871 150951
rect 215198 147737 218871 148023
rect 215198 147650 218864 147737
rect 215198 147003 216861 147650
rect 10765 128929 11213 128945
rect 33333 128937 33781 128941
rect 10765 128373 11238 128929
rect 10790 128357 11238 128373
rect 33320 128369 33781 128937
rect 10968 128307 11045 128357
rect 10968 128103 11046 128307
rect 13010 128203 13515 128368
rect 33320 128365 33768 128369
rect 11149 128183 13515 128203
rect 11149 128150 11157 128183
rect 11191 128150 13515 128183
rect 11149 128141 13515 128150
rect 10968 128028 10974 128103
rect 11038 128028 11046 128103
rect 10968 128019 11046 128028
rect 11076 128103 11154 128113
rect 11076 128028 11083 128103
rect 11147 128028 11154 128103
rect 11076 127916 11154 128028
rect 11075 127896 11154 127916
rect 11193 128103 11281 128114
rect 11193 128028 11199 128103
rect 11274 128028 11281 128103
rect 11193 128016 11281 128028
rect 11075 127839 11153 127896
rect 10873 127771 11153 127839
rect 11193 127853 11271 128016
rect 11193 127802 11691 127853
rect 10873 127763 11152 127771
rect 10208 127762 11152 127763
rect 8981 127728 11152 127762
rect 11194 127733 11691 127802
rect 8981 127504 10949 127728
rect 11074 127725 11152 127728
rect 8980 127321 10949 127504
rect 8980 127319 10224 127321
rect 8980 126250 9482 127319
rect 8980 124650 9485 126250
rect 11256 124753 11691 127733
rect 13010 126755 13515 128141
rect 33468 128307 33545 128365
rect 33468 128103 33546 128307
rect 35510 128203 36015 128368
rect 55817 128367 56265 128939
rect 33649 128183 36015 128203
rect 33649 128150 33657 128183
rect 33691 128150 36015 128183
rect 33649 128141 36015 128150
rect 33468 128028 33474 128103
rect 33538 128028 33546 128103
rect 33468 128019 33546 128028
rect 33576 128103 33654 128113
rect 33576 128028 33583 128103
rect 33647 128028 33654 128103
rect 33576 127916 33654 128028
rect 33696 128103 33784 128114
rect 33696 128028 33702 128103
rect 33777 128028 33784 128103
rect 33696 128018 33784 128028
rect 33575 127896 33654 127916
rect 33693 128016 33784 128018
rect 33575 127839 33653 127896
rect 33373 127771 33653 127839
rect 33693 127853 33771 128016
rect 33693 127802 34191 127853
rect 31479 127762 32255 127764
rect 33373 127763 33652 127771
rect 32708 127762 33652 127763
rect 31479 127728 33652 127762
rect 33694 127733 34191 127802
rect 31479 127321 33449 127728
rect 33574 127725 33652 127728
rect 31479 127319 32724 127321
rect 31479 126249 32255 127319
rect 11244 124181 11692 124753
rect 31480 124650 31985 126249
rect 33756 124870 34191 127733
rect 35510 126755 36015 128141
rect 55968 128307 56045 128367
rect 55968 128103 56046 128307
rect 58010 128204 58515 128368
rect 78291 128351 78739 128923
rect 57750 128203 58515 128204
rect 56149 128183 58515 128203
rect 56149 128150 56157 128183
rect 56191 128150 58515 128183
rect 56149 128141 58515 128150
rect 55968 128028 55974 128103
rect 56038 128028 56046 128103
rect 55968 128019 56046 128028
rect 56076 128103 56154 128113
rect 56076 128028 56083 128103
rect 56147 128028 56154 128103
rect 56076 127916 56154 128028
rect 56075 127896 56154 127916
rect 56203 128103 56291 128114
rect 56203 128028 56209 128103
rect 56284 128028 56291 128103
rect 56203 128016 56291 128028
rect 56075 127839 56153 127896
rect 55873 127771 56153 127839
rect 56203 127853 56281 128016
rect 56203 127802 56691 127853
rect 55873 127763 56152 127771
rect 55208 127762 56152 127763
rect 53983 127755 54481 127761
rect 54745 127755 56152 127762
rect 53983 127728 56152 127755
rect 56204 127733 56691 127802
rect 53983 127327 55949 127728
rect 56074 127725 56152 127728
rect 56225 127626 56691 127733
rect 53983 126250 54481 127327
rect 54745 127321 55949 127327
rect 54745 127319 55224 127321
rect 33756 124650 34207 124870
rect 53980 124650 54485 126250
rect 56256 124939 56691 127626
rect 58010 126755 58515 128141
rect 78468 128307 78545 128351
rect 78468 128103 78546 128307
rect 80510 128203 81015 128368
rect 100767 128361 101215 128946
rect 78649 128183 81015 128203
rect 78649 128150 78657 128183
rect 78691 128150 81015 128183
rect 78649 128141 81015 128150
rect 78468 128028 78474 128103
rect 78538 128028 78546 128103
rect 78468 128019 78546 128028
rect 78576 128103 78654 128113
rect 78576 128028 78583 128103
rect 78647 128028 78654 128103
rect 78576 127916 78654 128028
rect 78575 127896 78654 127916
rect 78728 128103 78816 128114
rect 78728 128028 78734 128103
rect 78809 128028 78816 128103
rect 78728 128016 78816 128028
rect 78575 127839 78653 127896
rect 78373 127771 78653 127839
rect 78728 127853 78806 128016
rect 78728 127802 79191 127853
rect 76480 127761 76989 127764
rect 78373 127763 78652 127771
rect 77708 127762 78652 127763
rect 77245 127761 78652 127762
rect 76480 127728 78652 127761
rect 78729 127733 79191 127802
rect 76480 127321 78449 127728
rect 78574 127725 78652 127728
rect 76480 127320 77724 127321
rect 56241 124767 56691 124939
rect 76480 126242 76989 127320
rect 77245 127319 77724 127320
rect 56240 124650 56696 124767
rect 76480 124650 76985 126242
rect 78756 124907 79191 127733
rect 80510 126755 81015 128141
rect 100968 128307 101045 128361
rect 100968 128103 101046 128307
rect 103010 128203 103515 128368
rect 123305 128360 123753 128932
rect 101149 128183 103515 128203
rect 101149 128150 101157 128183
rect 101191 128150 103515 128183
rect 101149 128141 103515 128150
rect 100968 128028 100974 128103
rect 101038 128028 101046 128103
rect 100968 128019 101046 128028
rect 101076 128103 101154 128113
rect 101076 128028 101083 128103
rect 101147 128028 101154 128103
rect 101278 128103 101366 128114
rect 101278 128031 101284 128103
rect 101076 127916 101154 128028
rect 101075 127896 101154 127916
rect 101277 128028 101284 128031
rect 101359 128028 101366 128103
rect 101277 128016 101366 128028
rect 101075 127839 101153 127896
rect 101277 127853 101357 128016
rect 100873 127771 101153 127839
rect 100873 127763 101152 127771
rect 100208 127762 101152 127763
rect 99745 127760 101152 127762
rect 99230 127750 101152 127760
rect 98977 127728 101152 127750
rect 101273 127732 101691 127853
rect 98977 127321 100949 127728
rect 101074 127725 101152 127728
rect 98977 126250 99481 127321
rect 99745 127319 100224 127321
rect 98977 126223 99485 126250
rect 78751 124815 79199 124907
rect 78744 124650 79199 124815
rect 98980 124650 99485 126223
rect 101256 124843 101691 127732
rect 103010 126755 103515 128141
rect 123468 128307 123545 128360
rect 123468 128103 123546 128307
rect 125510 128203 126015 128368
rect 145780 128345 146228 128917
rect 123649 128183 126015 128203
rect 123649 128150 123657 128183
rect 123649 128149 123691 128150
rect 123860 128149 126015 128183
rect 123649 128141 126015 128149
rect 125242 128140 126015 128141
rect 123468 128028 123474 128103
rect 123538 128028 123546 128103
rect 123468 128019 123546 128028
rect 123576 128103 123654 128113
rect 123576 128028 123583 128103
rect 123647 128028 123654 128103
rect 123576 127916 123654 128028
rect 123575 127896 123654 127916
rect 123878 128103 123966 128114
rect 123878 128028 123884 128103
rect 123959 128098 123966 128103
rect 123959 128028 123971 128098
rect 123575 127839 123653 127896
rect 123878 127853 123971 128028
rect 123373 127771 123653 127839
rect 123373 127763 123652 127771
rect 122708 127762 123652 127763
rect 121480 127728 123652 127762
rect 121480 127321 123449 127728
rect 123574 127725 123652 127728
rect 121480 127320 122724 127321
rect 101246 124781 101691 124843
rect 121480 126250 121960 127320
rect 122245 127319 122724 127320
rect 101246 124650 101699 124781
rect 121480 124650 121985 126250
rect 123756 124970 124191 127853
rect 125510 126755 126015 128140
rect 145968 128307 146045 128345
rect 145968 128103 146046 128307
rect 148010 128203 148515 128368
rect 168346 128354 168794 128926
rect 146149 128183 148515 128203
rect 146149 128150 146157 128183
rect 146149 128148 146178 128150
rect 146552 128148 148515 128183
rect 146149 128141 148515 128148
rect 145968 128028 145974 128103
rect 146038 128028 146046 128103
rect 145968 128019 146046 128028
rect 146076 128103 146154 128113
rect 146076 128028 146083 128103
rect 146147 128028 146154 128103
rect 146578 128103 146666 128114
rect 146578 128081 146584 128103
rect 146076 127916 146154 128028
rect 146075 127896 146154 127916
rect 146577 128028 146584 128081
rect 146659 128081 146666 128103
rect 146659 128028 146667 128081
rect 146075 127839 146153 127896
rect 146577 127853 146667 128028
rect 145873 127771 146153 127839
rect 145873 127763 146152 127771
rect 145208 127762 146152 127763
rect 143980 127728 146152 127762
rect 143980 127321 145949 127728
rect 146074 127725 146152 127728
rect 143980 127319 145224 127321
rect 143980 127318 144920 127319
rect 143980 126250 144484 127318
rect 123756 124846 124205 124970
rect 123738 124650 124205 124846
rect 143980 124650 144485 126250
rect 146256 124728 146691 127853
rect 148010 126755 148515 128141
rect 168468 128307 168545 128354
rect 168468 128103 168546 128307
rect 170510 128203 171015 128368
rect 189801 128354 190249 128926
rect 208375 128767 213588 129003
rect 208371 128543 213588 128767
rect 168649 128183 171015 128203
rect 168649 128150 168657 128183
rect 168649 128148 168680 128150
rect 169445 128148 171015 128183
rect 168649 128141 171015 128148
rect 168468 128028 168474 128103
rect 168538 128028 168546 128103
rect 168468 128019 168546 128028
rect 168576 128103 168654 128113
rect 168576 128028 168583 128103
rect 168647 128028 168654 128103
rect 168576 127916 168654 128028
rect 169478 128103 169566 128114
rect 169478 128028 169484 128103
rect 169559 128028 169566 128103
rect 169478 128016 169566 128028
rect 168575 127896 168654 127916
rect 169480 127896 169566 128016
rect 168575 127839 168653 127896
rect 168373 127771 168653 127839
rect 166480 127762 166985 127764
rect 168373 127763 168652 127771
rect 167708 127762 168652 127763
rect 166480 127728 168652 127762
rect 166480 127321 168449 127728
rect 168574 127725 168652 127728
rect 166480 127320 167724 127321
rect 33759 124298 34207 124650
rect 56241 124367 56689 124650
rect 78751 124335 79199 124650
rect 101251 124209 101699 124650
rect 123757 124398 124205 124650
rect 146255 124156 146703 124728
rect 166480 124650 166985 127320
rect 167245 127319 167724 127320
rect 169435 124931 169912 127896
rect 170510 126755 171015 128141
rect 189967 128120 190046 128354
rect 193010 128204 193515 128368
rect 208371 128367 208741 128543
rect 208371 128365 208710 128367
rect 208371 128204 208568 128365
rect 192749 128203 193515 128204
rect 190171 128184 193515 128203
rect 190171 128150 190186 128184
rect 192127 128150 193515 128184
rect 190171 128141 193515 128150
rect 190171 128137 192166 128141
rect 189968 128103 190046 128120
rect 189968 128028 189974 128103
rect 190038 128028 190046 128103
rect 189968 128019 190046 128028
rect 190076 128103 190154 128113
rect 190076 128028 190083 128103
rect 190147 128028 190154 128103
rect 192178 128103 192266 128114
rect 192178 128066 192184 128103
rect 190076 127916 190154 128028
rect 190075 127896 190154 127916
rect 192177 128028 192184 128066
rect 192259 128028 192266 128103
rect 190075 127869 190153 127896
rect 189429 127867 190153 127869
rect 188985 127734 190153 127867
rect 192177 127824 192266 128028
rect 192177 127797 192267 127824
rect 188985 126250 189484 127734
rect 190075 127733 190153 127734
rect 192178 127606 192267 127797
rect 192177 127555 192267 127606
rect 192177 127132 192266 127555
rect 192177 127107 192267 127132
rect 192178 126904 192267 127107
rect 169415 124650 169912 124931
rect 188980 124650 189485 126250
rect 192104 124846 192426 126904
rect 193010 126755 193515 128141
rect 208467 128136 208544 128204
rect 215510 128203 216015 128368
rect 213649 128200 216015 128203
rect 208668 128183 218657 128200
rect 208668 128178 213657 128183
rect 213691 128178 218657 128183
rect 208668 128148 208679 128178
rect 218645 128148 218657 128178
rect 208668 128138 218657 128148
rect 208467 128133 208546 128136
rect 208468 128103 208546 128133
rect 208468 128028 208474 128103
rect 208538 128028 208546 128103
rect 208468 128019 208546 128028
rect 208576 128103 208654 128113
rect 208576 128028 208583 128103
rect 208647 128028 208654 128103
rect 208576 127916 208654 128028
rect 208575 127896 208654 127916
rect 208575 127881 208653 127896
rect 208576 127865 208653 127881
rect 208524 126238 208750 127865
rect 215510 126755 216015 128138
rect 218678 128103 218766 128114
rect 218678 128099 218684 128103
rect 218677 128028 218684 128099
rect 218759 128028 218766 128103
rect 218677 127951 218766 128028
rect 211480 126238 211985 126250
rect 208524 125062 211985 126238
rect 208524 125056 208750 125062
rect 169415 124359 169863 124650
rect 192040 124274 192488 124846
rect 211480 124650 211985 125062
rect 218625 125023 218871 127951
rect 215896 125008 218871 125023
rect 215087 124737 218871 125008
rect 215087 124650 218864 124737
rect 215087 123986 216944 124650
rect 145717 105995 146147 106013
rect 10847 105337 11277 105977
rect 10968 105307 11045 105337
rect 10968 105103 11046 105307
rect 13010 105203 13515 105368
rect 33297 105342 33727 105982
rect 11149 105183 13515 105203
rect 11149 105150 11157 105183
rect 11191 105150 13515 105183
rect 11149 105141 13515 105150
rect 10968 104963 10974 105103
rect 11038 104963 11046 105103
rect 10968 104954 11046 104963
rect 11076 105103 11154 105113
rect 11076 104963 11083 105103
rect 11147 104963 11154 105103
rect 11076 104916 11154 104963
rect 11075 104896 11154 104916
rect 11193 105103 11281 105114
rect 11193 104963 11199 105103
rect 11274 104963 11281 105103
rect 11193 104951 11281 104963
rect 11075 104839 11153 104896
rect 10873 104771 11153 104839
rect 11193 104853 11271 104951
rect 11193 104802 11691 104853
rect 10873 104763 11152 104771
rect 10208 104762 11152 104763
rect 8981 104728 11152 104762
rect 11194 104733 11691 104802
rect 8981 104504 10949 104728
rect 11074 104725 11152 104728
rect 8980 104321 10949 104504
rect 8980 104319 10224 104321
rect 8980 103250 9482 104319
rect 8980 101650 9485 103250
rect 11256 101889 11691 104733
rect 13010 103755 13515 105141
rect 33468 105307 33545 105342
rect 33468 105103 33546 105307
rect 35510 105203 36015 105368
rect 55800 105352 56230 105992
rect 33649 105183 36015 105203
rect 33649 105150 33657 105183
rect 33691 105150 36015 105183
rect 33649 105141 36015 105150
rect 33468 104963 33474 105103
rect 33538 104963 33546 105103
rect 33468 104954 33546 104963
rect 33576 105103 33654 105113
rect 33576 104963 33583 105103
rect 33647 104963 33654 105103
rect 33696 105103 33784 105114
rect 33696 105018 33702 105103
rect 33576 104916 33654 104963
rect 33575 104896 33654 104916
rect 33693 104963 33702 105018
rect 33777 104963 33784 105103
rect 33693 104951 33784 104963
rect 33575 104839 33653 104896
rect 33373 104771 33653 104839
rect 33693 104853 33771 104951
rect 33693 104802 34191 104853
rect 31479 104762 32255 104764
rect 33373 104763 33652 104771
rect 32708 104762 33652 104763
rect 31479 104728 33652 104762
rect 33694 104733 34191 104802
rect 31479 104321 33449 104728
rect 33574 104725 33652 104728
rect 31479 104319 32724 104321
rect 31479 103249 32255 104319
rect 11256 101782 11956 101889
rect 11188 101249 11956 101782
rect 31480 101650 31985 103249
rect 33756 101910 34191 104733
rect 35510 103755 36015 105141
rect 55968 105307 56045 105352
rect 55968 105103 56046 105307
rect 58010 105204 58515 105368
rect 78289 105346 78719 105986
rect 57750 105203 58515 105204
rect 56149 105183 58515 105203
rect 56149 105150 56157 105183
rect 56191 105150 58515 105183
rect 56149 105141 58515 105150
rect 55968 104963 55974 105103
rect 56038 104963 56046 105103
rect 55968 104954 56046 104963
rect 56076 105103 56154 105113
rect 56076 104963 56083 105103
rect 56147 104963 56154 105103
rect 56076 104916 56154 104963
rect 56075 104896 56154 104916
rect 56203 105103 56291 105114
rect 56203 104963 56209 105103
rect 56284 104963 56291 105103
rect 56203 104951 56291 104963
rect 56075 104839 56153 104896
rect 55873 104771 56153 104839
rect 56203 104853 56281 104951
rect 56203 104802 56691 104853
rect 55873 104763 56152 104771
rect 55208 104762 56152 104763
rect 53983 104755 54481 104761
rect 54745 104755 56152 104762
rect 53983 104728 56152 104755
rect 56204 104733 56691 104802
rect 53983 104327 55949 104728
rect 56074 104725 56152 104728
rect 56225 104626 56691 104733
rect 53983 103250 54481 104327
rect 54745 104321 55949 104327
rect 54745 104319 55224 104321
rect 33756 101650 34203 101910
rect 53980 101650 54485 103250
rect 56256 101957 56691 104626
rect 58010 103755 58515 105141
rect 78468 105307 78545 105346
rect 78468 105103 78546 105307
rect 80510 105203 81015 105368
rect 100759 105355 101189 105995
rect 78649 105183 81015 105203
rect 78649 105150 78657 105183
rect 78691 105150 81015 105183
rect 78649 105141 81015 105150
rect 78468 104963 78474 105103
rect 78538 104963 78546 105103
rect 78468 104954 78546 104963
rect 78576 105103 78654 105113
rect 78576 104963 78583 105103
rect 78647 104963 78654 105103
rect 78576 104916 78654 104963
rect 78575 104896 78654 104916
rect 78728 105103 78816 105114
rect 78728 104963 78734 105103
rect 78809 104963 78816 105103
rect 78728 104951 78816 104963
rect 78575 104839 78653 104896
rect 78373 104771 78653 104839
rect 78728 104853 78806 104951
rect 78728 104802 79191 104853
rect 76480 104761 76989 104764
rect 78373 104763 78652 104771
rect 77708 104762 78652 104763
rect 77245 104761 78652 104762
rect 76480 104728 78652 104761
rect 78729 104733 79191 104802
rect 76480 104321 78449 104728
rect 78574 104725 78652 104728
rect 76480 104320 77724 104321
rect 76480 103242 76989 104320
rect 77245 104319 77724 104320
rect 56256 101767 56714 101957
rect 56240 101650 56714 101767
rect 76480 101650 76985 103242
rect 78756 101859 79191 104733
rect 80510 103755 81015 105141
rect 100968 105307 101045 105355
rect 100968 105103 101046 105307
rect 103010 105203 103515 105368
rect 123238 105346 123668 105986
rect 145708 105373 146147 105995
rect 101149 105183 103515 105203
rect 101149 105150 101157 105183
rect 101191 105150 103515 105183
rect 101149 105141 103515 105150
rect 100968 104963 100974 105103
rect 101038 104963 101046 105103
rect 100968 104954 101046 104963
rect 101076 105103 101154 105113
rect 101076 104963 101083 105103
rect 101147 104963 101154 105103
rect 101278 105103 101366 105114
rect 101278 105031 101284 105103
rect 101076 104916 101154 104963
rect 101075 104896 101154 104916
rect 101277 104963 101284 105031
rect 101359 104963 101366 105103
rect 101277 104951 101366 104963
rect 101075 104839 101153 104896
rect 101277 104853 101357 104951
rect 100873 104771 101153 104839
rect 100873 104763 101152 104771
rect 100208 104762 101152 104763
rect 99745 104760 101152 104762
rect 99230 104750 101152 104760
rect 98977 104728 101152 104750
rect 101273 104732 101691 104853
rect 98977 104321 100949 104728
rect 101074 104725 101152 104728
rect 98977 103250 99481 104321
rect 99745 104319 100224 104321
rect 98977 103223 99485 103250
rect 78756 101815 79196 101859
rect 78744 101650 79196 101815
rect 98980 101650 99485 103223
rect 101256 101843 101691 104732
rect 103010 103755 103515 105141
rect 123468 105307 123545 105346
rect 123468 105103 123546 105307
rect 125510 105203 126015 105368
rect 145708 105355 146138 105373
rect 123649 105183 126015 105203
rect 123649 105150 123657 105183
rect 123649 105149 123691 105150
rect 123860 105149 126015 105183
rect 123649 105141 126015 105149
rect 125242 105140 126015 105141
rect 123468 104963 123474 105103
rect 123538 104963 123546 105103
rect 123468 104954 123546 104963
rect 123576 105103 123654 105113
rect 123576 104963 123583 105103
rect 123647 104963 123654 105103
rect 123576 104916 123654 104963
rect 123575 104896 123654 104916
rect 123878 105103 123966 105114
rect 123878 104963 123884 105103
rect 123959 105098 123966 105103
rect 123959 104963 123971 105098
rect 123575 104839 123653 104896
rect 123878 104853 123971 104963
rect 123373 104771 123653 104839
rect 123373 104763 123652 104771
rect 122708 104762 123652 104763
rect 121480 104728 123652 104762
rect 121480 104321 123449 104728
rect 123574 104725 123652 104728
rect 121480 104320 122724 104321
rect 101246 101841 101691 101843
rect 101245 101650 101691 101841
rect 121480 103250 121960 104320
rect 122245 104319 122724 104320
rect 121480 101650 121985 103250
rect 123756 101846 124191 104853
rect 125510 103755 126015 105140
rect 145968 105307 146045 105355
rect 145968 105103 146046 105307
rect 148010 105203 148515 105368
rect 168268 105337 168698 105977
rect 146149 105183 148515 105203
rect 146149 105150 146157 105183
rect 146149 105148 146178 105150
rect 146552 105148 148515 105183
rect 146149 105141 148515 105148
rect 145968 104963 145974 105103
rect 146038 104963 146046 105103
rect 145968 104954 146046 104963
rect 146076 105103 146154 105113
rect 146076 104963 146083 105103
rect 146147 104963 146154 105103
rect 146578 105103 146666 105114
rect 146578 105081 146584 105103
rect 146076 104916 146154 104963
rect 146075 104896 146154 104916
rect 146577 104963 146584 105081
rect 146659 105081 146666 105103
rect 146659 104963 146667 105081
rect 146075 104839 146153 104896
rect 146577 104853 146667 104963
rect 145873 104771 146153 104839
rect 145873 104763 146152 104771
rect 145208 104762 146152 104763
rect 143980 104728 146152 104762
rect 143980 104321 145949 104728
rect 146074 104725 146152 104728
rect 143980 104319 145224 104321
rect 143980 104318 144920 104319
rect 143980 103250 144484 104318
rect 123738 101650 124200 101846
rect 143980 101650 144485 103250
rect 146256 101706 146691 104853
rect 148010 103755 148515 105141
rect 168468 105307 168545 105337
rect 168468 105103 168546 105307
rect 170510 105203 171015 105368
rect 189711 105346 190141 105986
rect 208262 105553 213037 106030
rect 168649 105183 171015 105203
rect 168649 105150 168657 105183
rect 168649 105148 168680 105150
rect 169445 105148 171015 105183
rect 168649 105141 171015 105148
rect 168468 104963 168474 105103
rect 168538 104963 168546 105103
rect 168468 104954 168546 104963
rect 168576 105103 168654 105113
rect 168576 104963 168583 105103
rect 168647 104963 168654 105103
rect 168576 104916 168654 104963
rect 169478 105103 169566 105114
rect 169478 104963 169484 105103
rect 169559 104963 169566 105103
rect 169478 104951 169566 104963
rect 168575 104896 168654 104916
rect 169480 104896 169566 104951
rect 168575 104839 168653 104896
rect 168373 104771 168653 104839
rect 166480 104762 166985 104764
rect 168373 104763 168652 104771
rect 167708 104762 168652 104763
rect 166480 104728 168652 104762
rect 166480 104321 168449 104728
rect 168574 104725 168652 104728
rect 166480 104320 167724 104321
rect 146221 101650 146691 101706
rect 166480 101650 166985 104320
rect 167245 104319 167724 104320
rect 169435 101904 169912 104896
rect 170510 103755 171015 105141
rect 189967 105120 190046 105346
rect 193010 105204 193515 105368
rect 208262 105355 208954 105553
rect 208371 105352 208954 105355
rect 208371 105204 208568 105352
rect 192749 105203 193515 105204
rect 190171 105184 193515 105203
rect 190171 105150 190186 105184
rect 192127 105150 193515 105184
rect 190171 105141 193515 105150
rect 190171 105137 192166 105141
rect 189968 105103 190046 105120
rect 189968 104963 189974 105103
rect 190038 104963 190046 105103
rect 189968 104954 190046 104963
rect 190076 105103 190154 105113
rect 190076 104963 190083 105103
rect 190147 104963 190154 105103
rect 192178 105103 192266 105114
rect 192178 105066 192184 105103
rect 190076 104916 190154 104963
rect 190075 104896 190154 104916
rect 192177 104963 192184 105066
rect 192259 104963 192266 105103
rect 190075 104869 190153 104896
rect 189429 104867 190153 104869
rect 188985 104734 190153 104867
rect 192177 104824 192266 104963
rect 192177 104797 192267 104824
rect 188985 103250 189484 104734
rect 190075 104733 190153 104734
rect 192178 104606 192267 104797
rect 192177 104555 192267 104606
rect 192177 104132 192266 104555
rect 192177 104107 192267 104132
rect 192178 103904 192267 104107
rect 169430 101650 169912 101904
rect 188980 101650 189485 103250
rect 192104 102021 192426 103904
rect 193010 103755 193515 105141
rect 208467 105136 208544 105204
rect 215510 105203 216015 105368
rect 213649 105200 216015 105203
rect 208668 105183 218657 105200
rect 208668 105178 213657 105183
rect 213691 105178 218657 105183
rect 208668 105148 208679 105178
rect 218645 105148 218657 105178
rect 208668 105138 218657 105148
rect 208467 105133 208546 105136
rect 208468 105103 208546 105133
rect 208468 104963 208474 105103
rect 208538 104963 208546 105103
rect 208468 104954 208546 104963
rect 208576 105103 208654 105113
rect 208576 104963 208583 105103
rect 208647 104963 208654 105103
rect 208576 104916 208654 104963
rect 208575 104896 208654 104916
rect 208575 104881 208653 104896
rect 208576 104865 208653 104881
rect 208524 103238 208750 104865
rect 215510 103755 216015 105138
rect 218678 105103 218766 105114
rect 218678 105099 218684 105103
rect 218677 104963 218684 105099
rect 218759 104963 218766 105103
rect 218677 104951 218766 104963
rect 211480 103238 211985 103250
rect 208524 102062 211985 103238
rect 208524 102056 208750 102062
rect 192104 101650 192537 102021
rect 211480 101650 211985 102062
rect 213956 102023 217235 102075
rect 218625 102023 218871 104951
rect 213956 101737 218871 102023
rect 213956 101650 218864 101737
rect 33773 101270 34203 101650
rect 56266 101317 56714 101650
rect 56266 101313 56696 101317
rect 11188 101142 11618 101249
rect 78766 101219 79196 101650
rect 101245 101201 101675 101650
rect 123742 101201 124172 101650
rect 146221 101066 146651 101650
rect 169430 101264 169860 101650
rect 192107 101381 192537 101650
rect 213956 100967 217235 101650
rect 10841 82349 11242 82670
rect 10968 82307 11045 82349
rect 10968 82103 11046 82307
rect 13010 82203 13515 82368
rect 33316 82344 33756 82899
rect 11149 82183 13515 82203
rect 11149 82150 11157 82183
rect 11191 82150 13515 82183
rect 11149 82141 13515 82150
rect 10968 81840 10974 82103
rect 11038 81840 11046 82103
rect 11076 82103 11154 82113
rect 11076 81916 11083 82103
rect 10970 81830 11045 81840
rect 11075 81828 11083 81916
rect 11147 81828 11154 82103
rect 11075 81816 11154 81828
rect 11193 82103 11281 82114
rect 11193 81828 11199 82103
rect 11274 81853 11281 82103
rect 11274 81828 11691 81853
rect 11075 81815 11153 81816
rect 10873 81771 11153 81815
rect 11193 81802 11691 81828
rect 10873 81763 11152 81771
rect 10208 81762 11152 81763
rect 8981 81728 11152 81762
rect 11194 81733 11691 81802
rect 8981 81504 10949 81728
rect 11074 81725 11152 81728
rect 8980 81321 10949 81504
rect 8980 81319 10224 81321
rect 8980 80250 9482 81319
rect 8980 78650 9485 80250
rect 11256 79022 11691 81733
rect 13010 80755 13515 82141
rect 33468 82307 33545 82344
rect 33468 82103 33546 82307
rect 35510 82203 36015 82368
rect 55807 82344 56247 82899
rect 33649 82183 36015 82203
rect 33649 82150 33657 82183
rect 33691 82150 36015 82183
rect 33649 82141 36015 82150
rect 33468 81845 33474 82103
rect 33538 81845 33546 82103
rect 33576 82103 33654 82113
rect 33576 81916 33583 82103
rect 33470 81830 33545 81845
rect 33575 81828 33583 81916
rect 33647 81828 33654 82103
rect 33696 82103 33784 82114
rect 33696 82018 33702 82103
rect 33575 81816 33654 81828
rect 33693 81828 33702 82018
rect 33777 81853 33784 82103
rect 33777 81828 34191 81853
rect 33575 81815 33653 81816
rect 33373 81771 33653 81815
rect 33693 81802 34191 81828
rect 31479 81762 32255 81764
rect 33373 81763 33652 81771
rect 32708 81762 33652 81763
rect 31479 81728 33652 81762
rect 33694 81733 34191 81802
rect 31479 81321 33449 81728
rect 33574 81725 33652 81728
rect 31479 81319 32724 81321
rect 31479 80249 32255 81319
rect 11238 78026 11705 79022
rect 31480 78650 31985 80249
rect 33756 79304 34191 81733
rect 35510 80755 36015 82141
rect 55968 82307 56045 82344
rect 55968 82103 56046 82307
rect 58010 82204 58515 82368
rect 78184 82344 78624 82899
rect 57750 82203 58515 82204
rect 56149 82183 58515 82203
rect 56149 82150 56157 82183
rect 56191 82150 58515 82183
rect 56149 82141 58515 82150
rect 55968 81845 55974 82103
rect 56038 81845 56046 82103
rect 56076 82103 56154 82113
rect 56076 81916 56083 82103
rect 55970 81830 56045 81845
rect 56075 81828 56083 81916
rect 56147 81828 56154 82103
rect 56075 81816 56154 81828
rect 56203 82103 56291 82114
rect 56203 81828 56209 82103
rect 56284 81853 56291 82103
rect 56284 81828 56691 81853
rect 56075 81815 56153 81816
rect 55873 81771 56153 81815
rect 56203 81802 56691 81828
rect 55873 81763 56152 81771
rect 55208 81762 56152 81763
rect 53983 81755 54481 81761
rect 54745 81755 56152 81762
rect 53983 81728 56152 81755
rect 56204 81733 56691 81802
rect 53983 81327 55949 81728
rect 56074 81725 56152 81728
rect 56225 81626 56691 81733
rect 53983 80250 54481 81327
rect 54745 81321 55949 81327
rect 54745 81319 55224 81321
rect 33756 78308 34223 79304
rect 53980 78650 54485 80250
rect 56256 78810 56691 81626
rect 58010 80755 58515 82141
rect 78468 82307 78545 82344
rect 78468 82103 78546 82307
rect 80510 82203 81015 82368
rect 100755 82362 101195 82917
rect 78649 82183 81015 82203
rect 78649 82150 78657 82183
rect 78691 82150 81015 82183
rect 78649 82141 81015 82150
rect 78468 81845 78474 82103
rect 78465 81840 78474 81845
rect 78538 81840 78546 82103
rect 78576 82103 78654 82113
rect 78576 81916 78583 82103
rect 78465 81825 78545 81840
rect 78575 81839 78583 81916
rect 78565 81828 78583 81839
rect 78647 81828 78654 82103
rect 78565 81816 78654 81828
rect 78728 82103 78816 82114
rect 78728 81828 78734 82103
rect 78809 81853 78816 82103
rect 78809 81828 79191 81853
rect 78565 81810 78653 81816
rect 78373 81771 78653 81810
rect 78728 81802 79191 81828
rect 76480 81761 76989 81764
rect 78373 81763 78652 81771
rect 77708 81762 78652 81763
rect 77245 81761 78652 81762
rect 76480 81728 78652 81761
rect 78729 81733 79191 81802
rect 76480 81321 78449 81728
rect 78574 81725 78652 81728
rect 76480 81320 77724 81321
rect 56213 78767 56691 78810
rect 76480 80242 76989 81320
rect 77245 81319 77724 81320
rect 56213 78650 56696 78767
rect 76480 78650 76985 80242
rect 78756 78871 79191 81733
rect 80510 80755 81015 82141
rect 100968 82307 101045 82362
rect 100968 82103 101046 82307
rect 103010 82203 103515 82368
rect 123273 82353 123713 82908
rect 101149 82183 103515 82203
rect 101149 82150 101157 82183
rect 101191 82150 103515 82183
rect 101149 82141 103515 82150
rect 100968 81840 100974 82103
rect 101038 81840 101046 82103
rect 101076 82103 101154 82113
rect 101076 81916 101083 82103
rect 100970 81830 101045 81840
rect 101075 81828 101083 81916
rect 101147 81828 101154 82103
rect 101278 82103 101366 82114
rect 101278 82031 101284 82103
rect 101277 81853 101284 82031
rect 101075 81816 101154 81828
rect 101273 81828 101284 81853
rect 101359 81853 101366 82103
rect 101359 81828 101691 81853
rect 101075 81815 101153 81816
rect 100873 81771 101153 81815
rect 100873 81763 101152 81771
rect 100208 81762 101152 81763
rect 99745 81760 101152 81762
rect 99230 81750 101152 81760
rect 98977 81728 101152 81750
rect 101273 81732 101691 81828
rect 98977 81321 100949 81728
rect 101074 81725 101152 81728
rect 98977 80250 99481 81321
rect 99745 81319 100224 81321
rect 98977 80223 99485 80250
rect 78740 78650 79191 78871
rect 98980 78650 99485 80223
rect 101256 78843 101691 81732
rect 103010 80755 103515 82141
rect 123468 82307 123545 82353
rect 123468 82103 123546 82307
rect 125510 82203 126015 82368
rect 145659 82344 146099 82899
rect 123649 82183 126015 82203
rect 123649 82150 123657 82183
rect 123649 82149 123691 82150
rect 123860 82149 126015 82183
rect 123649 82141 126015 82149
rect 125242 82140 126015 82141
rect 123468 81850 123474 82103
rect 123465 81845 123474 81850
rect 123538 81845 123546 82103
rect 123576 82103 123654 82113
rect 123576 81916 123583 82103
rect 123465 81830 123545 81845
rect 123575 81839 123583 81916
rect 123565 81828 123583 81839
rect 123647 81828 123654 82103
rect 123878 82103 123966 82114
rect 123878 81853 123884 82103
rect 123565 81816 123654 81828
rect 123756 81828 123884 81853
rect 123959 82098 123966 82103
rect 123959 81853 123971 82098
rect 123959 81828 124191 81853
rect 123565 81810 123653 81816
rect 123373 81771 123653 81810
rect 123373 81763 123652 81771
rect 122708 81762 123652 81763
rect 121480 81728 123652 81762
rect 121480 81321 123449 81728
rect 123574 81725 123652 81728
rect 121480 81320 122724 81321
rect 101246 78775 101691 78843
rect 101231 78650 101691 78775
rect 121480 80250 121960 81320
rect 122245 81319 122724 81320
rect 121480 78650 121985 80250
rect 123756 78846 124191 81828
rect 125510 80755 126015 82140
rect 145968 82307 146045 82344
rect 145968 82103 146046 82307
rect 148010 82203 148515 82368
rect 168327 82344 168767 82899
rect 189752 82882 190192 82943
rect 189744 82388 190192 82882
rect 207917 82556 212377 83499
rect 146149 82183 148515 82203
rect 146149 82150 146157 82183
rect 146149 82148 146178 82150
rect 146552 82148 148515 82183
rect 146149 82141 148515 82148
rect 145968 81845 145974 82103
rect 145965 81840 145974 81845
rect 146038 81840 146046 82103
rect 146076 82103 146154 82113
rect 146076 81916 146083 82103
rect 145965 81825 146045 81840
rect 146075 81828 146083 81916
rect 146147 81828 146154 82103
rect 146578 82103 146666 82114
rect 146578 82081 146584 82103
rect 146577 81853 146584 82081
rect 146075 81816 146154 81828
rect 146256 81828 146584 81853
rect 146659 82081 146666 82103
rect 146659 81853 146667 82081
rect 146659 81828 146691 81853
rect 146075 81800 146153 81816
rect 145873 81771 146153 81800
rect 145873 81763 146152 81771
rect 145208 81762 146152 81763
rect 143980 81728 146152 81762
rect 143980 81321 145949 81728
rect 146074 81725 146152 81728
rect 143980 81319 145224 81321
rect 143980 81318 144920 81319
rect 143980 80250 144484 81318
rect 123738 78819 124200 78846
rect 123738 78650 124216 78819
rect 143980 78650 144485 80250
rect 146256 78827 146691 81828
rect 148010 80755 148515 82141
rect 168468 82307 168545 82344
rect 168468 82103 168546 82307
rect 170510 82203 171015 82368
rect 189744 82327 190184 82388
rect 168649 82183 171015 82203
rect 168649 82150 168657 82183
rect 168649 82148 168680 82150
rect 169445 82148 171015 82183
rect 168649 82141 171015 82148
rect 168468 81845 168474 82103
rect 168538 81845 168546 82103
rect 168576 82103 168654 82113
rect 168576 81916 168583 82103
rect 168470 81825 168545 81845
rect 168575 81828 168583 81916
rect 168647 81828 168654 82103
rect 169478 82103 169566 82114
rect 169478 81896 169484 82103
rect 168575 81816 168654 81828
rect 169435 81828 169484 81896
rect 169559 81896 169566 82103
rect 169559 81828 169912 81896
rect 168575 81805 168653 81816
rect 168373 81771 168653 81805
rect 166480 81762 166985 81764
rect 168373 81763 168652 81771
rect 167708 81762 168652 81763
rect 166480 81728 168652 81762
rect 166480 81321 168449 81728
rect 168574 81725 168652 81728
rect 166480 81320 167724 81321
rect 146250 78650 146691 78827
rect 166480 78650 166985 81320
rect 167245 81319 167724 81320
rect 169435 78845 169912 81828
rect 170510 80755 171015 82141
rect 189967 82120 190046 82327
rect 193010 82204 193515 82368
rect 208357 82344 208710 82556
rect 208371 82204 208568 82344
rect 192749 82203 193515 82204
rect 190171 82184 193515 82203
rect 190171 82150 190186 82184
rect 192127 82150 193515 82184
rect 190171 82141 193515 82150
rect 190171 82137 192166 82141
rect 189968 82103 190046 82120
rect 189968 81880 189974 82103
rect 189965 81875 189974 81880
rect 190038 81875 190046 82103
rect 190076 82103 190154 82113
rect 190076 81916 190083 82103
rect 189429 81867 189940 81869
rect 188985 81800 189940 81867
rect 189965 81835 190045 81875
rect 190075 81828 190083 81916
rect 190147 81828 190154 82103
rect 192178 82103 192266 82114
rect 192178 82066 192184 82103
rect 190075 81816 190154 81828
rect 192177 81828 192184 82066
rect 192259 81828 192266 82103
rect 192177 81824 192266 81828
rect 190075 81800 190153 81816
rect 188985 81734 190153 81800
rect 192177 81797 192267 81824
rect 188985 80250 189484 81734
rect 190075 81733 190153 81734
rect 192178 81606 192267 81797
rect 192177 81555 192267 81606
rect 192177 81132 192266 81555
rect 192177 81107 192267 81132
rect 192178 80904 192267 81107
rect 169429 78650 169912 78845
rect 188980 78650 189485 80250
rect 192104 78995 192426 80904
rect 193010 80755 193515 82141
rect 208467 82136 208544 82204
rect 215510 82203 216015 82368
rect 213649 82200 216015 82203
rect 208668 82183 218657 82200
rect 208668 82178 213657 82183
rect 213691 82178 218657 82183
rect 208668 82148 208679 82178
rect 218645 82148 218657 82178
rect 208668 82138 218657 82148
rect 208467 82133 208546 82136
rect 208468 82103 208546 82133
rect 208468 81828 208474 82103
rect 208538 81865 208546 82103
rect 208576 82103 208654 82113
rect 208576 81916 208583 82103
rect 208575 81881 208583 81916
rect 208576 81865 208583 81881
rect 208538 81828 208545 81865
rect 208468 81820 208545 81828
rect 208580 81828 208583 81865
rect 208647 81865 208654 82103
rect 208647 81828 208750 81865
rect 208580 81785 208750 81828
rect 208524 80238 208750 81785
rect 215510 80755 216015 82138
rect 218678 82103 218766 82114
rect 218678 82099 218684 82103
rect 218677 81951 218684 82099
rect 218625 81828 218684 81951
rect 218759 81951 218766 82103
rect 218759 81828 218871 81951
rect 211480 80238 211985 80250
rect 208524 79062 211985 80238
rect 208524 79056 208750 79062
rect 56213 78255 56653 78650
rect 78740 78316 79180 78650
rect 101231 78220 101671 78650
rect 123776 78264 124216 78650
rect 146250 78272 146690 78650
rect 169429 78290 169869 78650
rect 192044 78440 192484 78995
rect 211480 78650 211985 79062
rect 218625 79023 218871 81828
rect 215896 78986 218871 79023
rect 214024 78737 218871 78986
rect 214024 78650 218864 78737
rect 214024 78043 218484 78650
rect 10876 59356 11238 59628
rect 10968 59307 11045 59356
rect 10968 59103 11046 59307
rect 13010 59203 13515 59368
rect 33313 59358 33748 59577
rect 11149 59183 13515 59203
rect 11149 59150 11157 59183
rect 11191 59150 13515 59183
rect 11149 59141 13515 59150
rect 10208 58762 10594 58763
rect 8981 58563 10594 58762
rect 10968 58633 10974 59103
rect 11038 58943 11046 59103
rect 11039 58633 11046 58943
rect 11076 59103 11154 59113
rect 11076 58941 11083 59103
rect 11147 58943 11154 59103
rect 10968 58627 11046 58633
rect 11078 58633 11083 58941
rect 11148 58941 11154 58943
rect 11193 59103 11281 59114
rect 11193 58941 11199 59103
rect 11274 58946 11281 59103
rect 11148 58633 11153 58941
rect 11078 58627 11153 58633
rect 11194 58633 11199 58941
rect 11275 58941 11281 58946
rect 11275 58889 11280 58941
rect 11275 58633 11694 58889
rect 11194 58628 11694 58633
rect 11079 58563 11153 58627
rect 8981 58504 11153 58563
rect 8980 58348 11153 58504
rect 8980 58321 11088 58348
rect 8980 58319 10224 58321
rect 10334 58319 11088 58321
rect 8980 57250 9482 58319
rect 11197 58148 11694 58628
rect 8980 55650 9485 57250
rect 11256 55973 11691 58148
rect 13010 57755 13515 59141
rect 33468 59307 33545 59358
rect 33468 59103 33546 59307
rect 35510 59203 36015 59368
rect 55667 59365 56218 59608
rect 33649 59183 36015 59203
rect 33649 59150 33657 59183
rect 33691 59150 36015 59183
rect 33649 59141 36015 59150
rect 31479 58762 32255 58764
rect 32708 58762 33120 58763
rect 31479 58592 33120 58762
rect 33468 58628 33474 59103
rect 33538 58628 33546 59103
rect 33576 59103 33654 59113
rect 33576 58916 33583 59103
rect 33575 58725 33583 58916
rect 33576 58683 33583 58725
rect 33468 58619 33546 58628
rect 33575 58628 33583 58683
rect 33647 58628 33654 59103
rect 33696 59103 33784 59114
rect 33696 59018 33702 59103
rect 33693 58802 33702 59018
rect 33694 58733 33702 58802
rect 33575 58592 33654 58628
rect 33696 58628 33702 58733
rect 33777 58853 33784 59103
rect 33777 58628 34191 58853
rect 33696 58616 34191 58628
rect 31479 58575 33654 58592
rect 31479 58334 33655 58575
rect 31479 58321 33595 58334
rect 31479 58319 32724 58321
rect 31479 57249 32255 58319
rect 11192 55405 11739 55973
rect 31480 55650 31985 57249
rect 33756 55882 34191 58616
rect 35510 57755 36015 59141
rect 55968 59307 56045 59365
rect 55968 59103 56046 59307
rect 58010 59204 58515 59368
rect 78358 59359 78746 59616
rect 57750 59203 58515 59204
rect 56149 59183 58515 59203
rect 56149 59150 56157 59183
rect 56191 59150 58515 59183
rect 56149 59141 58515 59150
rect 55208 58762 55657 58763
rect 53983 58755 54481 58761
rect 54745 58755 55657 58762
rect 53983 58560 55657 58755
rect 55968 58628 55974 59103
rect 56038 58628 56046 59103
rect 55968 58619 56046 58628
rect 56076 59103 56154 59113
rect 56076 58628 56083 59103
rect 56147 58628 56154 59103
rect 56076 58560 56154 58628
rect 56203 59103 56291 59114
rect 56203 58628 56209 59103
rect 56284 58997 56291 59103
rect 56284 58853 56568 58997
rect 56284 58628 56691 58853
rect 56203 58616 56691 58628
rect 53983 58327 56159 58560
rect 53983 57250 54481 58327
rect 54745 58321 56159 58327
rect 54745 58319 55224 58321
rect 55608 58317 56159 58321
rect 33689 55245 34273 55882
rect 53980 55650 54485 57250
rect 56256 55767 56691 58616
rect 58010 57755 58515 59141
rect 78468 59307 78545 59359
rect 78468 59103 78546 59307
rect 80510 59203 81015 59368
rect 100865 59352 101246 59639
rect 78649 59183 81015 59203
rect 78649 59150 78657 59183
rect 78691 59150 81015 59183
rect 78649 59141 81015 59150
rect 76480 58761 76989 58764
rect 77708 58762 78121 58763
rect 77245 58761 78121 58762
rect 76480 58557 78121 58761
rect 78468 58628 78474 59103
rect 78538 58628 78546 59103
rect 78576 59103 78654 59113
rect 78576 58916 78583 59103
rect 78575 58725 78583 58916
rect 78468 58619 78546 58628
rect 78576 58628 78583 58725
rect 78647 58628 78654 59103
rect 78576 58557 78654 58628
rect 78728 59103 78816 59114
rect 78728 58628 78734 59103
rect 78809 58992 78816 59103
rect 78809 58853 78980 58992
rect 78809 58628 79191 58853
rect 78728 58616 79191 58628
rect 76480 58321 78654 58557
rect 76480 58320 77724 58321
rect 76480 57242 76989 58320
rect 77245 58319 77724 58320
rect 56240 55669 56696 55767
rect 56186 55426 56737 55669
rect 76480 55650 76985 57242
rect 78756 55815 79191 58616
rect 80510 57755 81015 59141
rect 100968 59307 101045 59352
rect 100968 59103 101046 59307
rect 103010 59203 103515 59368
rect 123331 59353 123714 59685
rect 101149 59183 103515 59203
rect 101149 59150 101157 59183
rect 101191 59150 103515 59183
rect 101149 59141 103515 59150
rect 100208 58762 100539 58763
rect 99745 58760 100539 58762
rect 99230 58750 100539 58760
rect 98977 58561 100539 58750
rect 100968 58628 100974 59103
rect 101038 58628 101046 59103
rect 101076 59103 101154 59113
rect 101076 58916 101083 59103
rect 101075 58725 101083 58916
rect 100968 58619 101046 58628
rect 101076 58628 101083 58725
rect 101147 58628 101154 59103
rect 101278 59103 101366 59114
rect 101278 59031 101284 59103
rect 101277 58853 101284 59031
rect 101273 58732 101284 58853
rect 101076 58561 101154 58628
rect 98977 58509 101154 58561
rect 101256 58628 101284 58732
rect 101359 58853 101366 59103
rect 101359 58628 101691 58853
rect 98977 58321 101153 58509
rect 98977 57250 99481 58321
rect 99745 58319 100224 58321
rect 100509 58318 101153 58321
rect 98977 57223 99485 57250
rect 78744 55650 79191 55815
rect 98980 55650 99485 57223
rect 101256 56073 101691 58628
rect 103010 57755 103515 59141
rect 123468 59307 123545 59353
rect 123468 59103 123546 59307
rect 125510 59203 126015 59368
rect 145772 59361 146246 59789
rect 123649 59183 126015 59203
rect 123649 59150 123657 59183
rect 123649 59149 123691 59150
rect 123860 59149 126015 59183
rect 123649 59141 126015 59149
rect 125242 59140 126015 59141
rect 122708 58762 123196 58763
rect 121480 58561 123196 58762
rect 123468 58628 123474 59103
rect 123538 58628 123546 59103
rect 123576 59103 123654 59113
rect 123576 58916 123583 59103
rect 123575 58725 123583 58916
rect 123468 58619 123546 58628
rect 123576 58628 123583 58725
rect 123647 58628 123654 59103
rect 123878 59103 123966 59114
rect 123878 58853 123884 59103
rect 123576 58561 123654 58628
rect 121480 58478 123654 58561
rect 123877 58628 123884 58853
rect 123959 59098 123966 59103
rect 123959 58853 123971 59098
rect 123959 58628 124191 58853
rect 121480 58321 123651 58478
rect 121480 58320 122724 58321
rect 121480 57250 121960 58320
rect 122245 58319 122724 58320
rect 123039 58316 123651 58321
rect 123877 58115 124191 58628
rect 78746 55396 79191 55650
rect 101244 55298 101696 56073
rect 121480 55650 121985 57250
rect 123756 55912 124191 58115
rect 125510 57755 126015 59140
rect 145968 59307 146045 59361
rect 145968 59103 146046 59307
rect 148010 59203 148515 59368
rect 168139 59340 168843 60096
rect 146149 59183 148515 59203
rect 146149 59150 146157 59183
rect 146149 59148 146178 59150
rect 146552 59148 148515 59183
rect 146149 59141 148515 59148
rect 145208 58762 145562 58763
rect 143980 58541 145562 58762
rect 145968 58628 145974 59103
rect 146038 58628 146046 59103
rect 146076 59103 146154 59113
rect 146076 58916 146083 59103
rect 146075 58725 146083 58916
rect 145968 58619 146046 58628
rect 146076 58628 146083 58725
rect 146147 58628 146154 59103
rect 146578 59103 146666 59114
rect 146578 59081 146584 59103
rect 146076 58541 146154 58628
rect 143980 58525 146154 58541
rect 146577 58628 146584 59081
rect 146659 59081 146666 59103
rect 146659 58853 146667 59081
rect 146659 58628 146691 58853
rect 143980 58324 146151 58525
rect 143980 58321 145562 58324
rect 143980 58319 145224 58321
rect 143980 58318 144920 58319
rect 143980 57250 144484 58318
rect 146577 58044 146691 58628
rect 123581 55421 124385 55912
rect 143980 55650 144485 57250
rect 146256 55844 146691 58044
rect 148010 57755 148515 59141
rect 168468 59307 168545 59340
rect 168468 59103 168546 59307
rect 170510 59203 171015 59368
rect 189786 59355 191202 59651
rect 208343 59373 211752 60029
rect 168649 59183 171015 59203
rect 168649 59150 168657 59183
rect 168649 59148 168680 59150
rect 169445 59148 171015 59183
rect 168649 59141 171015 59148
rect 166480 58762 166985 58764
rect 167708 58762 168091 58763
rect 166480 58569 168091 58762
rect 168468 58628 168474 59103
rect 168538 58628 168546 59103
rect 168576 59103 168654 59113
rect 168576 58916 168583 59103
rect 168575 58725 168583 58916
rect 168468 58619 168546 58628
rect 168576 58628 168583 58725
rect 168647 58628 168654 59103
rect 169478 59103 169566 59114
rect 169478 58896 169484 59103
rect 168576 58569 168654 58628
rect 166480 58339 168654 58569
rect 169435 58628 169484 58896
rect 169559 58896 169566 59103
rect 169559 58628 169912 58896
rect 166480 58321 168649 58339
rect 166480 58320 167724 58321
rect 168066 58320 168649 58321
rect 146242 55416 146716 55844
rect 166480 55650 166985 58320
rect 167245 58319 167724 58320
rect 169435 55978 169912 58628
rect 170510 57755 171015 59141
rect 189967 59120 190046 59355
rect 193010 59204 193515 59368
rect 208352 59327 208757 59373
rect 208371 59204 208568 59327
rect 192749 59203 193515 59204
rect 190171 59184 193515 59203
rect 190171 59150 190186 59184
rect 192127 59150 193515 59184
rect 190171 59141 193515 59150
rect 190171 59137 192166 59141
rect 189968 59103 190046 59120
rect 189968 58628 189974 59103
rect 190038 58628 190046 59103
rect 190076 59103 190154 59113
rect 190076 58916 190083 59103
rect 189968 58619 190046 58628
rect 190075 58628 190083 58916
rect 190147 58628 190154 59103
rect 192178 59103 192266 59114
rect 192178 59066 192184 59103
rect 192177 58797 192184 59066
rect 190075 58616 190154 58628
rect 192178 58628 192184 58797
rect 192259 58824 192266 59103
rect 192259 58628 192267 58824
rect 190075 58530 190152 58616
rect 192178 58606 192267 58628
rect 188988 58417 190152 58530
rect 188985 58277 190152 58417
rect 192177 58555 192267 58606
rect 188985 58188 190150 58277
rect 188985 57250 189484 58188
rect 192177 58132 192266 58555
rect 192177 58107 192267 58132
rect 192178 57904 192267 58107
rect 169314 55222 170018 55978
rect 188980 55650 189485 57250
rect 192104 55767 192426 57904
rect 193010 57755 193515 59141
rect 208467 59136 208544 59204
rect 215510 59203 216015 59368
rect 213649 59200 216015 59203
rect 208668 59183 218657 59200
rect 208668 59178 213657 59183
rect 213691 59178 218657 59183
rect 208668 59148 208679 59178
rect 218645 59148 218657 59178
rect 208668 59138 218657 59148
rect 208467 59133 208546 59136
rect 208468 59103 208546 59133
rect 208468 58628 208474 59103
rect 208538 58865 208546 59103
rect 208576 59103 208654 59113
rect 208576 58916 208583 59103
rect 208575 58881 208583 58916
rect 208576 58865 208583 58881
rect 208538 58628 208547 58865
rect 208468 58619 208547 58628
rect 208524 58617 208547 58619
rect 208575 58628 208583 58865
rect 208647 58865 208654 59103
rect 208647 58628 208750 58865
rect 208575 58617 208750 58628
rect 208577 58562 208750 58617
rect 208524 57238 208750 58562
rect 215510 57755 216015 59138
rect 218678 59103 218766 59114
rect 218678 59099 218684 59103
rect 218677 58951 218684 59099
rect 218625 58628 218684 58951
rect 218759 58951 218766 59103
rect 218759 58628 218871 58951
rect 211480 57238 211985 57250
rect 208524 56062 211985 57238
rect 218625 56460 218871 58628
rect 208524 56056 208750 56062
rect 192061 55393 192447 55767
rect 211480 55650 211985 56062
rect 213788 55737 218871 56460
rect 213788 55650 218864 55737
rect 213788 55001 218839 55650
rect 10933 36344 11116 36607
rect 10968 36307 11045 36344
rect 10968 36103 11046 36307
rect 13010 36203 13515 36368
rect 33207 36342 33986 37065
rect 11149 36183 13515 36203
rect 11149 36150 11157 36183
rect 11191 36150 13515 36183
rect 11149 36141 13515 36150
rect 10968 35428 10974 36103
rect 11038 35428 11046 36103
rect 10968 35419 11046 35428
rect 11076 36103 11154 36113
rect 11076 35428 11083 36103
rect 11147 35428 11154 36103
rect 11076 35416 11154 35428
rect 11193 36103 11281 36114
rect 11193 35428 11199 36103
rect 11274 35814 11281 36103
rect 11274 35428 11695 35814
rect 11193 35416 11695 35428
rect 13010 35416 13515 36141
rect 33468 36307 33545 36342
rect 33468 36103 33546 36307
rect 35510 36203 36015 36368
rect 55837 36363 56211 36787
rect 33649 36183 36015 36203
rect 33649 36150 33657 36183
rect 33691 36150 36015 36183
rect 33649 36141 36015 36150
rect 33468 35428 33474 36103
rect 33538 35428 33546 36103
rect 33468 35419 33546 35428
rect 33576 36103 33654 36113
rect 33576 35428 33583 36103
rect 33647 35428 33654 36103
rect 33576 35416 33654 35428
rect 33696 36103 33784 36114
rect 33696 35428 33702 36103
rect 33777 35844 33784 36103
rect 33777 35830 33924 35844
rect 33777 35428 34112 35830
rect 33696 35416 34112 35428
rect 35510 35416 36015 36141
rect 55968 36307 56045 36363
rect 55968 36103 56046 36307
rect 58010 36204 58515 36368
rect 78194 36354 78691 36837
rect 57750 36203 58515 36204
rect 56149 36183 58515 36203
rect 56149 36150 56157 36183
rect 56191 36150 58515 36183
rect 56149 36141 58515 36150
rect 55968 35428 55974 36103
rect 56038 35428 56046 36103
rect 55968 35419 56046 35428
rect 56076 36103 56154 36113
rect 56076 35428 56083 36103
rect 56147 35428 56154 36103
rect 56076 35416 56154 35428
rect 56203 36103 56291 36114
rect 56203 35428 56209 36103
rect 56284 35865 56291 36103
rect 56284 35428 56618 35865
rect 56203 35416 56618 35428
rect 58010 35416 58515 36141
rect 78468 36307 78545 36354
rect 78468 36103 78546 36307
rect 80510 36203 81015 36368
rect 100777 36361 101214 36702
rect 78649 36183 81015 36203
rect 78649 36150 78657 36183
rect 78691 36150 81015 36183
rect 78649 36141 81015 36150
rect 78468 35428 78474 36103
rect 78538 35428 78546 36103
rect 78576 36103 78654 36113
rect 78576 35554 78583 36103
rect 78468 35419 78546 35428
rect 78575 35428 78583 35554
rect 78647 35428 78654 36103
rect 78575 35416 78654 35428
rect 78728 36103 78816 36114
rect 78728 35428 78734 36103
rect 78809 35757 78816 36103
rect 78809 35428 79001 35757
rect 78728 35416 79001 35428
rect 80510 35416 81015 36141
rect 100968 36307 101045 36361
rect 100968 36103 101046 36307
rect 103010 36203 103515 36368
rect 123260 36342 123795 37061
rect 101149 36183 103515 36203
rect 101149 36150 101157 36183
rect 101191 36150 103515 36183
rect 101149 36141 103515 36150
rect 100968 35428 100974 36103
rect 101038 35428 101046 36103
rect 100968 35419 101046 35428
rect 101076 36103 101154 36113
rect 101076 35428 101083 36103
rect 101147 35428 101154 36103
rect 101076 35416 101154 35428
rect 101278 36103 101366 36114
rect 101278 35428 101284 36103
rect 101359 35842 101366 36103
rect 101359 35428 101569 35842
rect 101278 35416 101569 35428
rect 103010 35416 103515 36141
rect 123468 36307 123545 36342
rect 123468 36103 123546 36307
rect 125510 36203 126015 36368
rect 145815 36356 146238 36779
rect 123649 36183 126015 36203
rect 123649 36150 123657 36183
rect 123649 36149 123691 36150
rect 123860 36149 126015 36183
rect 123649 36141 126015 36149
rect 125242 36140 126015 36141
rect 123468 35428 123474 36103
rect 123538 35428 123546 36103
rect 123576 36103 123654 36113
rect 123576 35605 123583 36103
rect 123468 35419 123546 35428
rect 123573 35428 123583 35605
rect 123647 35428 123654 36103
rect 123573 35416 123654 35428
rect 123878 36103 123966 36114
rect 123878 35428 123884 36103
rect 123959 36098 123966 36103
rect 123959 35741 123971 36098
rect 123959 35428 124041 35741
rect 123878 35416 124041 35428
rect 125510 35416 126015 36140
rect 145968 36307 146045 36356
rect 145968 36103 146046 36307
rect 148010 36203 148515 36368
rect 167870 36337 168739 36818
rect 146149 36183 148515 36203
rect 146149 36150 146157 36183
rect 146149 36148 146178 36150
rect 146552 36148 148515 36183
rect 146149 36141 148515 36148
rect 145968 35428 145974 36103
rect 146038 35428 146046 36103
rect 145968 35419 146046 35428
rect 146076 36103 146154 36113
rect 146076 35428 146083 36103
rect 146147 35428 146154 36103
rect 146076 35416 146154 35428
rect 146574 36103 146708 36114
rect 146574 35428 146584 36103
rect 146659 35946 146708 36103
rect 146659 35428 146737 35946
rect 11082 35299 11154 35416
rect 8981 35022 11154 35299
rect 8981 34732 11102 35022
rect 8980 34448 11102 34732
rect 8980 34250 9482 34448
rect 11207 34340 11695 35416
rect 33577 35193 33652 35416
rect 31525 35021 33652 35193
rect 31525 34732 33637 35021
rect 8980 32650 9485 34250
rect 11256 33013 11691 34340
rect 31479 34255 33637 34732
rect 33710 34732 34112 35416
rect 56084 35201 56141 35416
rect 53981 35083 56141 35201
rect 33710 34454 34191 34732
rect 53981 34470 56134 35083
rect 56225 34732 56618 35416
rect 78575 35039 78651 35416
rect 76485 34732 78651 35039
rect 78757 34732 79001 35416
rect 101081 35072 101147 35416
rect 98992 34998 101147 35072
rect 98992 34732 101136 34998
rect 101291 34732 101569 35416
rect 123573 35008 123651 35416
rect 121580 34732 123651 35008
rect 123890 34732 124041 35416
rect 146077 35011 146141 35416
rect 146574 35399 146737 35428
rect 148010 35416 148515 36141
rect 168468 36307 168545 36337
rect 168468 36103 168546 36307
rect 170510 36203 171015 36368
rect 189761 36315 190291 36584
rect 168649 36183 171015 36203
rect 168649 36150 168657 36183
rect 168649 36148 168680 36150
rect 169445 36148 171015 36183
rect 168649 36141 171015 36148
rect 168468 35428 168474 36103
rect 168538 35428 168546 36103
rect 168468 35419 168546 35428
rect 168576 36103 168654 36113
rect 168576 35428 168583 36103
rect 168647 35428 168654 36103
rect 168576 35416 168654 35428
rect 169478 36103 169566 36114
rect 169478 35428 169484 36103
rect 169559 35948 169566 36103
rect 169559 35428 169812 35948
rect 169478 35416 169812 35428
rect 170510 35416 171015 36141
rect 189967 36120 190046 36315
rect 193010 36204 193515 36368
rect 208354 36348 212665 36997
rect 208371 36204 208568 36348
rect 192749 36203 193515 36204
rect 190171 36184 193515 36203
rect 190171 36150 190186 36184
rect 192127 36150 193515 36184
rect 190171 36141 193515 36150
rect 190171 36137 192166 36141
rect 189968 36103 190046 36120
rect 189968 35428 189974 36103
rect 190038 35428 190046 36103
rect 189968 35419 190046 35428
rect 190076 36103 190154 36113
rect 190076 35428 190083 36103
rect 190147 35593 190154 36103
rect 192178 36103 192266 36114
rect 190147 35428 190159 35593
rect 190076 35416 190159 35428
rect 192178 35428 192184 36103
rect 192259 35973 192266 36103
rect 192259 35428 192426 35973
rect 192178 35416 192426 35428
rect 193010 35416 193515 36141
rect 208467 36136 208544 36204
rect 215510 36203 216015 36368
rect 213649 36200 216015 36203
rect 208668 36183 218657 36200
rect 208668 36178 213657 36183
rect 213691 36178 218657 36183
rect 208668 36148 208679 36178
rect 218645 36148 218657 36178
rect 208668 36138 218657 36148
rect 208467 36133 208546 36136
rect 208468 36103 208546 36133
rect 208468 35428 208474 36103
rect 208538 35428 208546 36103
rect 208468 35419 208546 35428
rect 208576 36103 208654 36113
rect 208576 35428 208583 36103
rect 208647 35428 208654 36103
rect 208576 35416 208654 35428
rect 215510 35416 216015 36138
rect 218676 36103 218766 36114
rect 218676 35428 218684 36103
rect 218759 36042 218766 36103
rect 218759 35428 219012 36042
rect 31479 34249 32255 34255
rect 11087 32290 11866 33013
rect 31480 32650 31985 34249
rect 33756 33104 34191 34454
rect 53983 34250 54481 34470
rect 56225 34426 56691 34732
rect 33720 32381 34499 33104
rect 53980 32650 54485 34250
rect 56256 33053 56691 34426
rect 76480 34645 78651 34732
rect 76480 34339 78634 34645
rect 76480 34242 76989 34339
rect 56172 32078 56822 33053
rect 76480 32650 76985 34242
rect 78756 33205 79191 34732
rect 98977 34613 101136 34732
rect 98977 34250 99481 34613
rect 98977 34223 99485 34250
rect 78639 32054 79419 33205
rect 98980 32650 99485 34223
rect 101256 33010 101691 34732
rect 101237 32650 101691 33010
rect 121480 34709 123651 34732
rect 121480 34237 123632 34709
rect 121480 32650 121985 34237
rect 123864 34171 124191 34732
rect 143962 34194 146141 35011
rect 146593 34732 146737 35399
rect 123756 32981 124191 34171
rect 123746 32846 124281 32981
rect 123738 32650 124281 32846
rect 143980 32650 144485 34194
rect 146568 34000 146737 34732
rect 166480 34728 166985 34732
rect 168576 34728 168646 35416
rect 169498 34732 169812 35416
rect 190078 35006 190159 35416
rect 166446 34191 168647 34728
rect 146568 33644 146691 34000
rect 146256 33060 146691 33644
rect 101237 32113 101683 32650
rect 123746 32262 124281 32650
rect 146238 32125 146716 33060
rect 166480 32650 166985 34191
rect 169435 33007 169912 34732
rect 188979 34345 190161 35006
rect 192203 34732 192426 35416
rect 208577 34732 208639 35416
rect 218676 35415 219012 35428
rect 218697 34732 219012 35415
rect 188985 34250 189484 34345
rect 169396 32650 169912 33007
rect 188980 32650 189485 34250
rect 192104 32917 192426 34732
rect 208524 34238 208750 34732
rect 211480 34238 211985 34250
rect 208524 33062 211985 34238
rect 208524 33056 208750 33062
rect 169396 32166 169905 32650
rect 192088 32126 192441 32917
rect 211480 32650 211985 33062
rect 218625 34005 219012 34732
rect 218625 33023 218871 34005
rect 215896 32978 218871 33023
rect 214645 32737 218871 32978
rect 214645 32650 218864 32737
rect 214645 31970 217758 32650
rect 10922 13424 11218 13816
rect 10921 13301 11219 13424
rect 10968 13103 11046 13301
rect 13010 13203 13515 13368
rect 33191 13342 33747 13743
rect 11149 13183 13515 13203
rect 11149 13150 11157 13183
rect 11191 13150 13515 13183
rect 11149 13141 13515 13150
rect 9172 10577 9928 11185
rect 9172 9840 10176 10577
rect 9217 9055 10176 9840
rect 9752 3030 10176 9055
rect 10968 3128 10974 13103
rect 11038 3128 11046 13103
rect 11076 13103 11154 13113
rect 11076 3138 11083 13103
rect 10968 3119 11046 3128
rect 11075 3128 11083 3138
rect 11147 3128 11154 13103
rect 11075 3116 11154 3128
rect 11193 13103 11281 13114
rect 11193 3128 11199 13103
rect 11274 3128 11281 13103
rect 13010 12719 13515 13141
rect 33468 13307 33545 13342
rect 33468 13103 33546 13307
rect 35510 13203 36015 13368
rect 55624 13329 56240 13843
rect 33649 13183 36015 13203
rect 33649 13150 33657 13183
rect 33691 13150 36015 13183
rect 33649 13141 36015 13150
rect 11193 3116 11281 3128
rect 11075 3030 11153 3116
rect 9752 2955 11153 3030
rect 31551 3026 31975 9781
rect 33468 3128 33474 13103
rect 33538 3128 33546 13103
rect 33468 3119 33546 3128
rect 33576 13103 33654 13113
rect 33576 3128 33583 13103
rect 33647 3128 33654 13103
rect 33576 3026 33654 3128
rect 33696 13103 33784 13114
rect 33696 3128 33702 13103
rect 33777 3128 33784 13103
rect 35510 12145 36015 13141
rect 55968 13103 56046 13329
rect 58010 13204 58515 13368
rect 77978 13353 78742 13800
rect 57750 13203 58515 13204
rect 56149 13183 58515 13203
rect 56149 13150 56157 13183
rect 56191 13150 58515 13183
rect 56149 13141 58515 13150
rect 33696 3116 33784 3128
rect 31551 2996 33654 3026
rect 53915 3032 54493 10407
rect 55968 3128 55974 13103
rect 56038 3128 56046 13103
rect 55968 3119 56046 3128
rect 56076 13103 56154 13113
rect 56076 3128 56083 13103
rect 56147 3128 56154 13103
rect 56076 3032 56154 3128
rect 56203 13103 56291 13114
rect 56203 3128 56209 13103
rect 56284 3128 56291 13103
rect 58010 12539 58515 13141
rect 78468 13307 78545 13353
rect 78468 13103 78546 13307
rect 80510 13203 81015 13368
rect 100593 13341 101248 13949
rect 78649 13183 81015 13203
rect 78649 13150 78657 13183
rect 78691 13150 81015 13183
rect 78649 13141 81015 13150
rect 56203 3116 56291 3128
rect 76608 3078 76986 10846
rect 78468 3128 78474 13103
rect 78538 3128 78546 13103
rect 78468 3119 78546 3128
rect 78576 13103 78654 13113
rect 78576 3128 78583 13103
rect 78647 3128 78654 13103
rect 78576 3078 78654 3128
rect 78728 13103 78816 13114
rect 78728 3128 78734 13103
rect 78809 3128 78816 13103
rect 80510 12585 81015 13141
rect 100968 13307 101045 13341
rect 100968 13103 101046 13307
rect 103010 13203 103515 13368
rect 122926 13359 123745 13810
rect 101149 13183 103515 13203
rect 101149 13150 101157 13183
rect 101191 13150 103515 13183
rect 101149 13141 103515 13150
rect 78728 3116 78816 3128
rect 9752 2755 11146 2955
rect 9867 2753 11146 2755
rect 31551 2665 33648 2996
rect 53915 2661 56156 3032
rect 76608 3009 78654 3078
rect 98931 3028 99491 10748
rect 100968 3128 100974 13103
rect 101038 3128 101046 13103
rect 100968 3119 101046 3128
rect 101076 13103 101154 13113
rect 101076 3128 101083 13103
rect 101147 3128 101154 13103
rect 101076 3028 101154 3128
rect 101278 13103 101366 13114
rect 101278 3128 101284 13103
rect 101359 3128 101366 13103
rect 103010 12713 103515 13141
rect 123468 13307 123545 13359
rect 123468 13103 123546 13307
rect 125510 13203 126015 13368
rect 145461 13361 146244 13652
rect 123649 13183 126015 13203
rect 123649 13150 123657 13183
rect 123649 13149 123691 13150
rect 123860 13149 126015 13183
rect 123649 13141 126015 13149
rect 125242 13140 126015 13141
rect 101278 3116 101366 3128
rect 76608 2644 78651 3009
rect 98931 2608 101154 3028
rect 121419 3037 121964 10751
rect 123468 3128 123474 13103
rect 123538 3128 123546 13103
rect 123468 3119 123546 3128
rect 123576 13103 123654 13113
rect 123576 3128 123583 13103
rect 123647 3128 123654 13103
rect 123576 3037 123654 3128
rect 123878 13103 123966 13114
rect 123878 3128 123884 13103
rect 123959 13098 123966 13103
rect 123959 13077 123971 13098
rect 123959 3128 124014 13077
rect 125510 12199 126015 13140
rect 145968 13307 146045 13361
rect 145968 13103 146046 13307
rect 148010 13203 148515 13368
rect 167914 13359 168718 13880
rect 146149 13183 148515 13203
rect 146149 13150 146157 13183
rect 146149 13148 146178 13150
rect 146552 13148 148515 13183
rect 146149 13141 148515 13148
rect 146578 13113 146666 13114
rect 123878 3116 124014 3128
rect 123931 3082 124014 3116
rect 121419 2979 123654 3037
rect 143922 3072 144486 10752
rect 145968 3128 145974 13103
rect 146038 3128 146046 13103
rect 145968 3119 146046 3128
rect 146076 13103 146154 13113
rect 146076 3128 146083 13103
rect 146147 3128 146154 13103
rect 146076 3072 146154 3128
rect 121419 2592 123650 2979
rect 143922 2974 146154 3072
rect 146564 13103 146691 13113
rect 146564 3128 146584 13103
rect 146659 3128 146691 13103
rect 148010 12577 148515 13141
rect 168468 13307 168545 13359
rect 168468 13103 168546 13307
rect 170510 13203 171015 13368
rect 189802 13361 190873 13959
rect 168649 13183 171015 13203
rect 168649 13150 168657 13183
rect 168649 13148 168680 13150
rect 169445 13148 171015 13183
rect 168649 13141 171015 13148
rect 146564 3040 146691 3128
rect 166453 3038 167005 10655
rect 168468 3128 168474 13103
rect 168538 3128 168546 13103
rect 168468 3119 168546 3128
rect 168576 13103 168654 13113
rect 168576 3128 168583 13103
rect 168647 3128 168654 13103
rect 168576 3038 168654 3128
rect 169478 13103 169566 13114
rect 169478 3128 169484 13103
rect 169559 3128 169566 13103
rect 170510 12469 171015 13141
rect 189967 13120 190046 13361
rect 193010 13204 193515 13368
rect 208370 13361 212740 14128
rect 208371 13204 208568 13361
rect 192749 13203 193515 13204
rect 190171 13184 193515 13203
rect 190171 13150 190186 13184
rect 192127 13150 193515 13184
rect 190171 13141 193515 13150
rect 190171 13137 192166 13141
rect 189968 13103 190046 13120
rect 169478 3116 169566 3128
rect 143922 2641 146149 2974
rect 166453 2950 168654 3038
rect 188939 3044 189507 10879
rect 189968 3128 189974 13103
rect 190038 3128 190046 13103
rect 189968 3119 190046 3128
rect 190076 13103 190154 13113
rect 190076 3128 190083 13103
rect 190147 3128 190154 13103
rect 190076 3116 190154 3128
rect 192178 13103 192266 13114
rect 192178 3128 192184 13103
rect 192259 3128 192266 13103
rect 193010 12390 193515 13141
rect 208467 13136 208544 13204
rect 215510 13203 216015 13368
rect 213649 13200 216015 13203
rect 208668 13183 218657 13200
rect 208668 13178 213657 13183
rect 213691 13178 218657 13183
rect 208668 13148 208679 13178
rect 218645 13148 218657 13178
rect 208668 13138 218657 13148
rect 208467 13133 208546 13136
rect 208468 13103 208546 13133
rect 192178 3116 192266 3128
rect 193010 3116 193515 9510
rect 208468 3128 208474 13103
rect 208538 3128 208546 13103
rect 208468 3119 208546 3128
rect 208576 13103 208654 13113
rect 208576 3128 208583 13103
rect 208647 10167 208654 13103
rect 215510 12280 216015 13138
rect 218680 13111 218766 13114
rect 218680 13103 218894 13111
rect 218680 12947 218684 13103
rect 208647 8726 212418 10167
rect 218202 9939 218684 12947
rect 208647 3128 208654 8726
rect 215346 8527 218684 9939
rect 208576 3116 208654 3128
rect 218202 3128 218684 8527
rect 218759 3128 218894 13103
rect 190077 3044 190154 3116
rect 166453 2812 168652 2950
rect 188939 2897 190154 3044
rect 218202 2909 218894 3128
rect 188939 2678 190152 2897
<< metal5 >>
rect 22245 193650 22745 197368
rect 44745 193650 45245 197368
rect 67245 193650 67745 197368
rect 89745 193650 90245 197368
rect 112245 193650 112745 197368
rect 134745 193650 135245 197368
rect 157245 193650 157745 197368
rect 179745 193650 180245 197368
rect 202245 193650 202745 197368
rect 22245 170650 22745 174368
rect 44745 170650 45245 174368
rect 67245 170650 67745 174368
rect 89745 170650 90245 174368
rect 112245 170650 112745 174368
rect 134745 170650 135245 174368
rect 157245 170650 157745 174368
rect 179745 170650 180245 174368
rect 202245 170650 202745 174368
rect 22245 147650 22745 151368
rect 44745 147650 45245 151368
rect 67245 147650 67745 151368
rect 89745 147650 90245 151368
rect 112245 147650 112745 151368
rect 134745 147650 135245 151368
rect 157245 147650 157745 151368
rect 179745 147650 180245 151368
rect 202245 147650 202745 151368
rect 22245 124650 22745 128368
rect 44745 124650 45245 128368
rect 67245 124650 67745 128368
rect 89745 124650 90245 128368
rect 112245 124650 112745 128368
rect 134745 124650 135245 128368
rect 157245 124650 157745 128368
rect 179745 124650 180245 128368
rect 202245 124650 202745 128368
rect 22245 101650 22745 105368
rect 44745 101650 45245 105368
rect 67245 101650 67745 105368
rect 89745 101650 90245 105368
rect 112245 101650 112745 105368
rect 134745 101650 135245 105368
rect 157245 101650 157745 105368
rect 179745 101650 180245 105368
rect 202245 101650 202745 105368
rect 22245 78650 22745 82368
rect 44745 78650 45245 82368
rect 67245 78650 67745 82368
rect 89745 78650 90245 82368
rect 112245 78650 112745 82368
rect 134745 78650 135245 82368
rect 157245 78650 157745 82368
rect 179745 78650 180245 82368
rect 202245 78650 202745 82368
rect 22245 55650 22745 59368
rect 44745 55650 45245 59368
rect 67245 55650 67745 59368
rect 89745 55650 90245 59368
rect 112245 55650 112745 59368
rect 134745 55650 135245 59368
rect 157245 55650 157745 59368
rect 179745 55650 180245 59368
rect 202245 55650 202745 59368
rect 22245 32650 22745 36368
rect 44745 32650 45245 36368
rect 67245 32650 67745 36368
rect 89745 32650 90245 36368
rect 112245 32650 112745 36368
rect 134745 32650 135245 36368
rect 157245 32650 157745 36368
rect 179745 32650 180245 36368
rect 202245 32650 202745 36368
rect 22245 3116 22745 13368
rect 44745 3116 45245 13368
rect 67245 3116 67745 13368
rect 89745 3116 90245 13368
rect 112245 3116 112745 13368
rect 134745 3116 135245 13368
rect 157245 3116 157745 13368
rect 179745 3116 180245 13368
rect 202245 3116 202745 13368
use BarePadArray10x10  BarePadArray10x10_0
timestamp 1663665281
transform 1 0 0 0 1 0
box -5 0 224995 230000
<< end >>
