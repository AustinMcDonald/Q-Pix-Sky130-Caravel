magic
tech sky130A
magscale 1 2
timestamp 1663455834
<< nwell >>
rect 4463 -2020 4910 -2017
rect -3870 -3340 4910 -2020
rect -3870 -4330 -1700 -3340
rect 2200 -3480 4910 -3340
rect 4463 -3482 4910 -3480
rect -1450 -6010 1290 -4690
<< pwell >>
rect -980 -4360 820 -3650
rect 3400 -4530 3810 -4480
rect 2210 -6010 4630 -4530
<< pmoslvt >>
rect -3400 -2790 -3330 -2190
rect -3400 -4260 -3330 -3060
rect -3130 -4260 -3060 -3060
rect -2860 -4260 -2790 -3060
rect -2590 -4260 -2520 -3060
rect -2320 -4260 -2250 -3060
rect -990 -3280 -920 -2080
rect -720 -3280 -650 -2080
rect -450 -3280 -380 -2080
rect 220 -3280 290 -2080
rect 490 -3280 560 -2080
rect 760 -3280 830 -2080
rect 2670 -3410 2740 -2210
rect 2940 -3410 3010 -2210
rect 3210 -3410 3280 -2210
rect 3480 -3410 3550 -2210
rect 3750 -3410 3820 -2210
rect 4020 -3410 4090 -2210
rect 4290 -3410 4360 -2210
rect -990 -5950 -920 -4750
rect -720 -5950 -650 -4750
rect -450 -5950 -380 -4750
rect 220 -5950 290 -4750
rect 490 -5950 560 -4750
rect 760 -5950 830 -4750
<< nmoslvt >>
rect -520 -4290 -450 -3690
rect -250 -4290 -180 -3690
rect 20 -4290 90 -3690
rect 290 -4290 360 -3690
rect 3760 -5870 3830 -4670
rect 4030 -5870 4100 -4670
rect 4300 -5870 4370 -4670
<< ndiff >>
rect -720 -3730 -520 -3690
rect -720 -4250 -700 -3730
rect -540 -4250 -520 -3730
rect -720 -4290 -520 -4250
rect -450 -3730 -250 -3690
rect -450 -4250 -430 -3730
rect -270 -4250 -250 -3730
rect -450 -4290 -250 -4250
rect -180 -3730 20 -3690
rect -180 -4250 -160 -3730
rect 0 -4250 20 -3730
rect -180 -4290 20 -4250
rect 90 -3730 290 -3690
rect 90 -4250 110 -3730
rect 270 -4250 290 -3730
rect 90 -4290 290 -4250
rect 360 -3730 560 -3690
rect 360 -4250 380 -3730
rect 540 -4250 560 -3730
rect 360 -4290 560 -4250
rect 3560 -4700 3760 -4670
rect 3560 -5830 3580 -4700
rect 3740 -5830 3760 -4700
rect 3560 -5870 3760 -5830
rect 3830 -4710 4030 -4670
rect 3830 -5330 3850 -4710
rect 4010 -4840 4030 -4710
rect 3830 -5830 3851 -5330
rect 4011 -5830 4030 -4840
rect 3830 -5870 4030 -5830
rect 4100 -4720 4300 -4670
rect 4100 -5830 4120 -4720
rect 4280 -5830 4300 -4720
rect 4100 -5870 4300 -5830
rect 4370 -4710 4570 -4670
rect 4370 -5330 4390 -4710
rect 4550 -4781 4570 -4710
rect 4370 -5831 4391 -5330
rect 4551 -5831 4570 -4781
rect 4370 -5870 4570 -5831
<< pdiff >>
rect -1190 -2120 -990 -2080
rect -3600 -2221 -3400 -2190
rect -3600 -2760 -3580 -2221
rect -3430 -2760 -3400 -2221
rect -3600 -2790 -3400 -2760
rect -3330 -2220 -2730 -2190
rect -3330 -2760 -3300 -2220
rect -2760 -2760 -2730 -2220
rect -3330 -2790 -2730 -2760
rect -3600 -3100 -3400 -3060
rect -3600 -4230 -3580 -3100
rect -3430 -4230 -3400 -3100
rect -3600 -4260 -3400 -4230
rect -3330 -3106 -3130 -3060
rect -3330 -3110 -3309 -3106
rect -3330 -4230 -3310 -3110
rect -3330 -4233 -3309 -4230
rect -3157 -4233 -3130 -3106
rect -3330 -4260 -3130 -4233
rect -3060 -3110 -2860 -3060
rect -3060 -4230 -3040 -3110
rect -2890 -4230 -2860 -3110
rect -3060 -4260 -2860 -4230
rect -2790 -3105 -2590 -3060
rect -2790 -4232 -2770 -3105
rect -2618 -4232 -2590 -3105
rect -2790 -4260 -2590 -4232
rect -2520 -3110 -2320 -3060
rect -2520 -4230 -2500 -3110
rect -2350 -4230 -2320 -3110
rect -2520 -4260 -2320 -4230
rect -2250 -3100 -2050 -3060
rect -2250 -4230 -2230 -3100
rect -2080 -4230 -2050 -3100
rect -2250 -4260 -2050 -4230
rect -1190 -3250 -1140 -2120
rect -1010 -3250 -990 -2120
rect -1190 -3280 -990 -3250
rect -920 -2120 -720 -2080
rect -920 -3250 -880 -2120
rect -750 -3250 -720 -2120
rect -920 -3280 -720 -3250
rect -650 -2120 -450 -2080
rect -650 -3250 -610 -2120
rect -480 -3250 -450 -2120
rect -650 -3280 -450 -3250
rect -380 -2120 -180 -2080
rect -380 -3250 -360 -2120
rect -230 -3250 -180 -2120
rect 20 -2120 220 -2080
rect -380 -3280 -180 -3250
rect 20 -3250 60 -2120
rect 190 -3250 220 -2120
rect 20 -3280 220 -3250
rect 290 -2120 490 -2080
rect 290 -3250 320 -2120
rect 450 -3250 490 -2120
rect 290 -3280 490 -3250
rect 560 -2110 760 -2080
rect 560 -3240 590 -2110
rect 720 -3240 760 -2110
rect 560 -3280 760 -3240
rect 830 -2110 1030 -2080
rect 830 -3240 850 -2110
rect 980 -3240 1030 -2110
rect 830 -3280 1030 -3240
rect 2470 -2250 2670 -2210
rect 2470 -3367 2490 -2250
rect 2650 -3000 2670 -2250
rect 2649 -3367 2670 -3000
rect 2470 -3410 2670 -3367
rect 2740 -2279 2940 -2210
rect 2740 -3385 2758 -2279
rect 2916 -2590 2940 -2279
rect 2740 -3390 2760 -3385
rect 2920 -3390 2940 -2590
rect 2740 -3410 2940 -3390
rect 3010 -2250 3210 -2210
rect 3010 -3000 3030 -2250
rect 3190 -2277 3210 -2250
rect 3010 -3384 3034 -3000
rect 3195 -3383 3210 -2277
rect 3193 -3384 3210 -3383
rect 3010 -3410 3210 -3384
rect 3280 -2246 3480 -2210
rect 3280 -3390 3300 -2246
rect 3459 -2590 3480 -2246
rect 3460 -3390 3480 -2590
rect 3280 -3393 3301 -3390
rect 3457 -3393 3480 -3390
rect 3280 -3410 3480 -3393
rect 3550 -2250 3750 -2210
rect 3550 -2287 3570 -2250
rect 3550 -3393 3569 -2287
rect 3730 -3000 3750 -2250
rect 3550 -3395 3570 -3393
rect 3729 -3395 3750 -3000
rect 3550 -3397 3572 -3395
rect 3728 -3397 3750 -3395
rect 3550 -3410 3750 -3397
rect 3820 -2257 4020 -2210
rect 3820 -2675 3839 -2257
rect 3998 -2282 4020 -2257
rect 3999 -2590 4020 -2282
rect 3820 -3038 3840 -2675
rect 3820 -3390 3838 -3038
rect 4000 -3390 4020 -2590
rect 3820 -3410 4020 -3390
rect 4090 -2250 4290 -2210
rect 4090 -3000 4110 -2250
rect 4270 -2277 4290 -2250
rect 4272 -2976 4290 -2277
rect 4090 -3383 4114 -3000
rect 4090 -3394 4115 -3383
rect 4090 -3397 4118 -3394
rect 4274 -3397 4290 -2976
rect 4090 -3410 4290 -3397
rect 4360 -2277 4560 -2210
rect 4360 -3390 4380 -2277
rect 4539 -2279 4560 -2277
rect 4540 -3390 4560 -2279
rect 4360 -3410 4560 -3390
rect -1190 -4790 -990 -4750
rect -1190 -5920 -1140 -4790
rect -1010 -5920 -990 -4790
rect -1190 -5950 -990 -5920
rect -920 -4790 -720 -4750
rect -920 -5920 -880 -4790
rect -750 -5920 -720 -4790
rect -920 -5950 -720 -5920
rect -650 -4790 -450 -4750
rect -650 -5920 -610 -4790
rect -480 -5920 -450 -4790
rect -650 -5950 -450 -5920
rect -380 -4790 -180 -4750
rect -380 -5920 -360 -4790
rect -230 -5920 -180 -4790
rect 20 -4790 220 -4750
rect -380 -5950 -180 -5920
rect 20 -5920 60 -4790
rect 190 -5920 220 -4790
rect 20 -5950 220 -5920
rect 290 -4790 490 -4750
rect 290 -5920 320 -4790
rect 450 -5920 490 -4790
rect 290 -5950 490 -5920
rect 560 -4780 760 -4750
rect 560 -5910 590 -4780
rect 720 -5910 760 -4780
rect 560 -5950 760 -5910
rect 830 -4780 1030 -4750
rect 830 -5910 850 -4780
rect 980 -5910 1030 -4780
rect 830 -5950 1030 -5910
<< ndiffc >>
rect -700 -4250 -540 -3730
rect -430 -4250 -270 -3730
rect -160 -4250 0 -3730
rect 110 -4250 270 -3730
rect 380 -4250 540 -3730
rect 3580 -5830 3740 -4700
rect 3850 -4840 4010 -4710
rect 3850 -5330 4011 -4840
rect 3851 -5830 4011 -5330
rect 4120 -5830 4280 -4720
rect 4390 -4781 4550 -4710
rect 4390 -5330 4551 -4781
rect 4391 -5831 4551 -5330
<< pdiffc >>
rect -3580 -2760 -3430 -2221
rect -3300 -2760 -2760 -2220
rect -3580 -4230 -3430 -3100
rect -3309 -3110 -3157 -3106
rect -3310 -4230 -3157 -3110
rect -3309 -4233 -3157 -4230
rect -3040 -4230 -2890 -3110
rect -2770 -4232 -2618 -3105
rect -2500 -4230 -2350 -3110
rect -2230 -4230 -2080 -3100
rect -1140 -3250 -1010 -2120
rect -880 -3250 -750 -2120
rect -610 -3250 -480 -2120
rect -360 -3250 -230 -2120
rect 60 -3250 190 -2120
rect 320 -3250 450 -2120
rect 590 -3240 720 -2110
rect 850 -3240 980 -2110
rect 2490 -3000 2650 -2250
rect 2490 -3367 2649 -3000
rect 2758 -2590 2916 -2279
rect 2758 -3385 2920 -2590
rect 2760 -3390 2920 -3385
rect 3030 -2277 3190 -2250
rect 3030 -3000 3195 -2277
rect 3034 -3383 3195 -3000
rect 3034 -3384 3193 -3383
rect 3300 -2590 3459 -2246
rect 3300 -3390 3460 -2590
rect 3301 -3393 3457 -3390
rect 3570 -2287 3730 -2250
rect 3569 -3000 3730 -2287
rect 3569 -3393 3729 -3000
rect 3570 -3395 3729 -3393
rect 3572 -3397 3728 -3395
rect 3839 -2282 3998 -2257
rect 3839 -2590 3999 -2282
rect 3839 -2675 4000 -2590
rect 3840 -3038 4000 -2675
rect 3838 -3390 4000 -3038
rect 4110 -2277 4270 -2250
rect 4110 -2976 4272 -2277
rect 4110 -3000 4274 -2976
rect 4114 -3383 4274 -3000
rect 4115 -3394 4274 -3383
rect 4118 -3397 4274 -3394
rect 4380 -2279 4539 -2277
rect 4380 -3390 4540 -2279
rect -1140 -5920 -1010 -4790
rect -880 -5920 -750 -4790
rect -610 -5920 -480 -4790
rect -360 -5920 -230 -4790
rect 60 -5920 190 -4790
rect 320 -5920 450 -4790
rect 590 -5910 720 -4780
rect 850 -5910 980 -4780
<< psubdiff >>
rect -920 -3730 -720 -3690
rect -920 -4250 -900 -3730
rect -740 -4250 -720 -3730
rect -920 -4290 -720 -4250
rect 560 -3730 760 -3690
rect 560 -4250 590 -3730
rect 750 -4250 760 -3730
rect 560 -4290 760 -4250
rect 3360 -4700 3560 -4670
rect 2900 -5150 3020 -5120
rect 2900 -5400 2930 -5150
rect 2990 -5400 3020 -5150
rect 2900 -5430 3020 -5400
rect 3360 -5830 3380 -4700
rect 3540 -5830 3560 -4700
rect 3360 -5870 3560 -5830
<< nsubdiff >>
rect -1390 -2120 -1190 -2080
rect -3800 -2221 -3600 -2190
rect -3800 -2760 -3780 -2221
rect -3630 -2760 -3600 -2221
rect -3800 -2790 -3600 -2760
rect -3800 -3100 -3600 -3060
rect -3800 -4230 -3780 -3100
rect -3630 -4230 -3600 -3100
rect -3800 -4260 -3600 -4230
rect -2050 -3092 -1750 -3060
rect -2050 -4236 -1959 -3092
rect -1795 -3552 -1750 -3092
rect -1390 -3250 -1360 -2120
rect -1230 -3250 -1190 -2120
rect -1390 -3280 -1190 -3250
rect -180 -2140 20 -2080
rect -180 -3240 -130 -2140
rect -30 -3240 20 -2140
rect -180 -3280 20 -3240
rect 1030 -2086 1230 -2080
rect 1030 -2110 1231 -2086
rect 1030 -3250 1080 -2110
rect 1210 -3250 1231 -2110
rect 1030 -3253 1231 -3250
rect 2270 -2250 2470 -2210
rect 2270 -2410 2290 -2250
rect 2440 -2410 2470 -2250
rect 2270 -3220 2291 -2410
rect 2438 -3220 2470 -2410
rect 1030 -3280 1230 -3253
rect 2270 -3380 2290 -3220
rect 2440 -3380 2470 -3220
rect 2270 -3410 2470 -3380
rect 4660 -2250 4860 -2210
rect 4660 -2410 4680 -2250
rect 4660 -3369 4682 -2410
rect 4832 -3369 4860 -2250
rect 4660 -3410 4860 -3369
rect -1795 -3693 -1745 -3552
rect -1795 -4236 -1746 -3693
rect -2050 -4250 -1746 -4236
rect -2050 -4260 -1750 -4250
rect -1390 -4790 -1190 -4750
rect -1390 -5920 -1360 -4790
rect -1230 -5920 -1190 -4790
rect -1390 -5950 -1190 -5920
rect -180 -4810 20 -4750
rect -180 -5910 -130 -4810
rect -30 -5910 20 -4810
rect -180 -5950 20 -5910
rect 1030 -4780 1230 -4750
rect 1030 -5920 1080 -4780
rect 1210 -5920 1230 -4780
rect 1030 -5950 1230 -5920
<< psubdiffcont >>
rect -900 -4250 -740 -3730
rect 590 -4250 750 -3730
rect 2930 -5400 2990 -5150
rect 3380 -5830 3540 -4700
<< nsubdiffcont >>
rect -3780 -2760 -3630 -2221
rect -3780 -4230 -3630 -3100
rect -1959 -4236 -1795 -3092
rect -1360 -3250 -1230 -2120
rect -130 -3240 -30 -2140
rect 1080 -3250 1210 -2110
rect 2290 -2410 2440 -2250
rect 2291 -3220 2438 -2410
rect 2290 -3380 2440 -3220
rect 4680 -2410 4832 -2250
rect 4682 -3369 4832 -2410
rect -1360 -5920 -1230 -4790
rect -130 -5910 -30 -4810
rect 1080 -5920 1210 -4780
<< poly >>
rect -990 -1900 -380 -1880
rect -990 -2000 -970 -1900
rect -400 -2000 -380 -1900
rect -990 -2020 -380 -2000
rect -990 -2080 -920 -2020
rect -720 -2080 -650 -2020
rect -450 -2080 -380 -2020
rect 220 -1900 830 -1880
rect 220 -2000 240 -1900
rect 810 -2000 830 -1900
rect 220 -2020 830 -2000
rect 220 -2080 290 -2020
rect 490 -2080 560 -2020
rect 760 -2080 830 -2020
rect 2670 -2040 4360 -2020
rect -3400 -2190 -3330 -2160
rect -3400 -2870 -3330 -2790
rect -3400 -2890 -2250 -2870
rect -3400 -2980 -3300 -2890
rect -2760 -2980 -2250 -2890
rect -3400 -3000 -2250 -2980
rect -3400 -3060 -3330 -3000
rect -3130 -3060 -3060 -3000
rect -2860 -3060 -2790 -3000
rect -2590 -3060 -2520 -3000
rect -2320 -3060 -2250 -3000
rect 2670 -2130 2690 -2040
rect 4340 -2130 4360 -2040
rect 2670 -2150 4360 -2130
rect 2670 -2210 2740 -2150
rect 2940 -2210 3010 -2150
rect 3210 -2210 3280 -2150
rect 3480 -2210 3550 -2150
rect 3750 -2210 3820 -2150
rect 4020 -2210 4090 -2150
rect 4290 -2210 4360 -2150
rect -990 -3340 -920 -3280
rect -720 -3340 -650 -3280
rect -450 -3340 -380 -3280
rect 220 -3340 290 -3280
rect 490 -3340 560 -3280
rect 760 -3340 830 -3280
rect 2670 -3450 2740 -3410
rect 2940 -3450 3010 -3410
rect 3210 -3450 3280 -3410
rect 3480 -3450 3550 -3410
rect 3750 -3450 3820 -3410
rect 4020 -3450 4090 -3410
rect 4290 -3450 4360 -3410
rect -520 -3560 360 -3530
rect -520 -3640 -430 -3560
rect -10 -3640 360 -3560
rect -520 -3650 360 -3640
rect -520 -3690 -450 -3650
rect -250 -3690 -180 -3650
rect 20 -3690 90 -3650
rect 290 -3690 360 -3650
rect -3400 -4300 -3330 -4260
rect -3130 -4300 -3060 -4260
rect -2860 -4300 -2790 -4260
rect -2590 -4300 -2520 -4260
rect -2320 -4300 -2250 -4260
rect -520 -4360 -450 -4290
rect -250 -4360 -180 -4290
rect 20 -4360 90 -4290
rect 290 -4360 360 -4290
rect -520 -4390 760 -4360
rect -520 -4480 380 -4390
rect 350 -4520 380 -4480
rect 730 -4520 760 -4390
rect 350 -4540 760 -4520
rect 3370 -4480 4370 -4470
rect -990 -4750 -920 -4690
rect -720 -4750 -650 -4690
rect -450 -4750 -380 -4690
rect 220 -4750 290 -4690
rect 490 -4750 560 -4690
rect 760 -4750 830 -4690
rect 3370 -4590 3400 -4480
rect 3810 -4490 4370 -4480
rect 4350 -4590 4370 -4490
rect 3370 -4610 4370 -4590
rect 3760 -4670 3830 -4610
rect 4030 -4670 4100 -4610
rect 4300 -4670 4370 -4610
rect -990 -6180 -920 -5950
rect -720 -6180 -650 -5950
rect -450 -6180 -380 -5950
rect 220 -6010 290 -5950
rect 490 -6010 560 -5950
rect 760 -6010 830 -5950
rect 3760 -5970 3830 -5870
rect 4030 -5970 4100 -5870
rect 4300 -5970 4370 -5870
rect 220 -6030 830 -6010
rect 220 -6130 240 -6030
rect 810 -6130 830 -6030
rect 220 -6150 830 -6130
rect -990 -6200 -380 -6180
rect -990 -6300 -970 -6200
rect -400 -6300 -380 -6200
rect -990 -6320 -380 -6300
<< polycont >>
rect -970 -2000 -400 -1900
rect 240 -2000 810 -1900
rect -3300 -2980 -2760 -2890
rect 2690 -2130 4340 -2040
rect -430 -3640 -10 -3560
rect 380 -4520 730 -4390
rect 3400 -4490 3810 -4480
rect 3400 -4590 4350 -4490
rect 240 -6130 810 -6030
rect -970 -6300 -400 -6200
<< xpolycontact >>
rect 2320 -5070 2720 -4560
rect 2320 -5980 2720 -5470
<< ppolyres >>
rect 2320 -5470 2720 -5070
<< locali >>
rect -990 -1900 -380 -1880
rect -990 -2000 -970 -1900
rect -400 -2000 -380 -1900
rect -990 -2020 -380 -2000
rect 220 -1900 830 -1880
rect 220 -2000 240 -1900
rect 810 -2000 830 -1900
rect 220 -2020 830 -2000
rect 2670 -2040 4360 -2020
rect -1390 -2120 -1210 -2090
rect -3801 -2221 -3418 -2191
rect -3801 -2593 -3780 -2221
rect -3800 -2760 -3780 -2593
rect -3630 -2760 -3580 -2221
rect -3430 -2403 -3418 -2221
rect -3320 -2220 -2740 -2200
rect -3430 -2760 -3420 -2403
rect -3800 -2780 -3420 -2760
rect -3320 -2760 -3300 -2220
rect -2760 -2760 -2740 -2220
rect -3320 -2890 -2740 -2760
rect -3320 -2980 -3300 -2890
rect -2760 -2980 -2740 -2890
rect -3320 -3000 -2740 -2980
rect -3800 -3100 -3430 -3080
rect -2790 -3090 -2591 -3087
rect -3800 -4230 -3780 -3100
rect -3630 -4230 -3580 -3100
rect -3330 -3106 -3130 -3090
rect -3330 -3110 -3309 -3106
rect -3330 -3610 -3310 -3110
rect -3800 -4250 -3430 -4230
rect -3329 -4230 -3310 -3610
rect -3329 -4233 -3309 -4230
rect -3157 -4233 -3130 -3106
rect -3060 -3110 -2860 -3090
rect -3060 -3111 -3040 -3110
rect -2890 -3111 -2860 -3110
rect -3060 -3610 -3041 -3111
rect -3059 -3710 -3041 -3610
rect -3329 -4250 -3130 -4233
rect -3060 -4234 -3041 -3710
rect -2889 -4234 -2860 -3111
rect -3060 -4250 -2860 -4234
rect -2790 -3105 -2590 -3090
rect -2790 -4232 -2770 -3105
rect -2618 -4232 -2590 -3105
rect -2520 -3091 -2320 -3090
rect -2520 -3109 -2318 -3091
rect -2520 -3610 -2504 -3109
rect -2352 -3110 -2318 -3109
rect -2519 -3710 -2504 -3610
rect -2790 -4250 -2590 -4232
rect -2520 -4232 -2504 -3710
rect -2350 -4230 -2318 -3110
rect -2250 -3100 -2050 -3080
rect -2250 -3101 -2230 -3100
rect -2250 -3610 -2234 -3101
rect -2352 -4232 -2318 -4230
rect -2520 -4250 -2318 -4232
rect -2249 -4228 -2234 -3610
rect -2249 -4230 -2230 -4228
rect -2080 -4230 -2050 -3100
rect -1978 -3092 -1771 -3075
rect -1978 -3691 -1959 -3092
rect -2249 -4250 -2050 -4230
rect -2790 -4252 -2591 -4250
rect -2518 -4254 -2318 -4250
rect -2248 -4256 -2050 -4250
rect -1982 -4236 -1959 -3691
rect -1795 -4236 -1771 -3092
rect -1390 -3250 -1360 -2120
rect -1230 -3250 -1210 -2120
rect -1390 -3270 -1210 -3250
rect -1170 -2120 -990 -2090
rect -1170 -3250 -1140 -2120
rect -1010 -3250 -990 -2120
rect -1170 -3270 -990 -3250
rect -910 -2120 -730 -2090
rect -910 -3250 -880 -2120
rect -750 -3250 -730 -2120
rect -910 -3270 -730 -3250
rect -640 -2120 -460 -2090
rect -640 -3250 -610 -2120
rect -480 -3250 -460 -2120
rect -640 -3270 -460 -3250
rect -380 -2120 -200 -2090
rect -380 -3250 -360 -2120
rect -230 -3250 -200 -2120
rect -380 -3270 -200 -3250
rect -150 -2140 -10 -2110
rect -150 -3240 -130 -2140
rect -30 -3240 -10 -2140
rect -150 -3260 -10 -3240
rect 40 -2120 220 -2090
rect 40 -3250 60 -2120
rect 190 -3250 220 -2120
rect 40 -3270 220 -3250
rect 300 -2120 480 -2090
rect 300 -3250 320 -2120
rect 450 -3250 480 -2120
rect 300 -3270 480 -3250
rect 570 -2110 750 -2090
rect 570 -3240 590 -2110
rect 720 -3240 750 -2110
rect 570 -3270 750 -3240
rect 830 -2110 1010 -2090
rect 830 -3240 850 -2110
rect 980 -3240 1010 -2110
rect 830 -3270 1010 -3240
rect 1050 -2110 1230 -2090
rect 1050 -3250 1080 -2110
rect 1210 -3250 1230 -2110
rect 2670 -2130 2690 -2040
rect 4340 -2130 4360 -2040
rect 2670 -2150 4360 -2130
rect 2276 -2216 2472 -2214
rect 2276 -2219 2667 -2216
rect 2276 -2230 2671 -2219
rect 2270 -2250 2671 -2230
rect 2270 -2410 2290 -2250
rect 2440 -2410 2490 -2250
rect 2270 -2430 2291 -2410
rect 2276 -3200 2291 -2430
rect 1050 -3270 1230 -3250
rect 2270 -3220 2291 -3200
rect 2438 -3220 2490 -2410
rect 2270 -3380 2290 -3220
rect 2440 -3367 2490 -3220
rect 2650 -3000 2671 -2250
rect 2742 -2279 2938 -2215
rect 2742 -2560 2758 -2279
rect 2649 -3367 2671 -3000
rect 2440 -3380 2671 -3367
rect 2270 -3400 2671 -3380
rect 2276 -3407 2671 -3400
rect 2464 -3409 2671 -3407
rect 2475 -3412 2671 -3409
rect 2740 -3385 2758 -2560
rect 2916 -2560 2938 -2279
rect 3007 -2230 3203 -2213
rect 3007 -2250 3210 -2230
rect 2916 -2590 2940 -2560
rect 2740 -3390 2760 -3385
rect 2920 -3390 2940 -2590
rect 2740 -3410 2940 -3390
rect 3007 -3000 3030 -2250
rect 3190 -2277 3210 -2250
rect 3007 -3384 3034 -3000
rect 3195 -3060 3210 -2277
rect 3281 -2246 3477 -2221
rect 3552 -2230 3748 -2217
rect 3281 -2560 3300 -2246
rect 3195 -3383 3203 -3060
rect 3193 -3384 3203 -3383
rect 3007 -3406 3203 -3384
rect 3280 -3390 3300 -2560
rect 3459 -2560 3477 -2246
rect 3550 -2250 3750 -2230
rect 3550 -2287 3570 -2250
rect 3459 -2590 3480 -2560
rect 3280 -3393 3301 -3390
rect 3460 -3390 3480 -2590
rect 3550 -3060 3569 -2287
rect 3730 -3000 3750 -2250
rect 3821 -2257 4017 -2216
rect 4091 -2230 4287 -2219
rect 3821 -2560 3839 -2257
rect 3998 -2282 4017 -2257
rect 3457 -3393 3480 -3390
rect 3280 -3410 3480 -3393
rect 3552 -3393 3569 -3060
rect 3552 -3395 3570 -3393
rect 3552 -3397 3572 -3395
rect 3729 -3060 3750 -3000
rect 3820 -2675 3839 -2560
rect 3820 -3038 3840 -2675
rect 3999 -2560 4017 -2282
rect 4090 -2250 4290 -2230
rect 3999 -2590 4020 -2560
rect 3729 -3395 3748 -3060
rect 3728 -3397 3748 -3395
rect 3552 -3410 3748 -3397
rect 3820 -3390 3838 -3038
rect 4000 -3390 4020 -2590
rect 4090 -3000 4110 -2250
rect 4270 -2277 4290 -2250
rect 4090 -3050 4114 -3000
rect 4272 -2976 4290 -2277
rect 4363 -2277 4559 -2211
rect 4363 -2560 4380 -2277
rect 4539 -2279 4559 -2277
rect 3820 -3410 4020 -3390
rect 4091 -3383 4114 -3050
rect 4274 -3050 4290 -2976
rect 4091 -3394 4115 -3383
rect 4091 -3397 4118 -3394
rect 4274 -3369 4287 -3050
rect 4274 -3397 4290 -3369
rect 3281 -3414 3477 -3410
rect 4091 -3412 4290 -3397
rect 4360 -3390 4380 -2560
rect 4540 -2560 4559 -2279
rect 4660 -2250 4860 -2230
rect 4660 -2410 4680 -2250
rect 4660 -2430 4682 -2410
rect 4540 -3390 4560 -2560
rect 4360 -3410 4560 -3390
rect 4663 -3369 4682 -2430
rect 4832 -3369 4860 -2250
rect 4663 -3406 4860 -3369
rect 4252 -3413 4290 -3412
rect -440 -3560 10 -3530
rect -440 -3640 -430 -3560
rect -10 -3640 10 -3560
rect -440 -3650 10 -3640
rect -1982 -4256 -1771 -4236
rect -920 -3730 -530 -3710
rect -920 -4250 -900 -3730
rect -740 -4250 -700 -3730
rect -540 -4250 -530 -3730
rect -920 -4270 -530 -4250
rect -440 -3730 -260 -3650
rect -440 -4250 -430 -3730
rect -270 -4250 -260 -3730
rect -440 -4270 -260 -4250
rect -170 -3730 10 -3710
rect -170 -4250 -160 -3730
rect 0 -4250 10 -3730
rect -170 -4270 10 -4250
rect 100 -3730 280 -3710
rect 100 -4250 110 -3730
rect 270 -4250 280 -3730
rect 100 -4270 280 -4250
rect 370 -3730 760 -3710
rect 370 -4250 380 -3730
rect 540 -4250 590 -3730
rect 750 -4250 760 -3730
rect 2100 -4020 2990 -3980
rect 2100 -4170 2370 -4020
rect 370 -4270 760 -4250
rect 350 -4390 760 -4360
rect 350 -4520 380 -4390
rect 730 -4520 760 -4390
rect 350 -4540 760 -4520
rect 2320 -4560 2370 -4170
rect 2960 -4420 2990 -4020
rect 2960 -4440 4370 -4420
rect 3670 -4480 4370 -4440
rect 3810 -4490 4370 -4480
rect 4350 -4590 4370 -4490
rect 3670 -4600 4370 -4590
rect -1390 -4790 -1210 -4760
rect -1390 -5920 -1360 -4790
rect -1230 -5920 -1210 -4790
rect -1390 -5940 -1210 -5920
rect -1170 -4790 -990 -4760
rect -1170 -5920 -1140 -4790
rect -1010 -5920 -990 -4790
rect -1170 -5940 -990 -5920
rect -910 -4790 -730 -4760
rect -910 -5920 -880 -4790
rect -750 -5920 -730 -4790
rect -910 -5940 -730 -5920
rect -640 -4790 -460 -4760
rect -640 -5920 -610 -4790
rect -480 -5920 -460 -4790
rect -640 -5940 -460 -5920
rect -380 -4790 -200 -4760
rect -380 -5920 -360 -4790
rect -230 -5920 -200 -4790
rect -380 -5940 -200 -5920
rect -150 -4810 -10 -4780
rect -150 -5910 -130 -4810
rect -30 -5910 -10 -4810
rect -150 -5930 -10 -5910
rect 40 -4790 220 -4760
rect 40 -5920 60 -4790
rect 190 -5920 220 -4790
rect 40 -5940 220 -5920
rect 300 -4790 480 -4760
rect 300 -5920 320 -4790
rect 450 -5920 480 -4790
rect 300 -5940 480 -5920
rect 570 -4780 750 -4760
rect 570 -5910 590 -4780
rect 720 -5910 750 -4780
rect 570 -5940 750 -5910
rect 830 -4780 1010 -4760
rect 830 -5910 850 -4780
rect 980 -5910 1010 -4780
rect 830 -5940 1010 -5910
rect 1050 -4780 1230 -4760
rect 1050 -5920 1080 -4780
rect 1210 -5920 1230 -4780
rect 2720 -4610 4370 -4600
rect 3532 -4680 3603 -4679
rect 3360 -4700 3760 -4680
rect 2910 -5150 3010 -5130
rect 2910 -5400 2930 -5150
rect 2990 -5400 3010 -5150
rect 2910 -5420 3010 -5400
rect 1050 -5940 1230 -5920
rect 3360 -5830 3380 -4700
rect 3540 -5830 3580 -4700
rect 3740 -5830 3760 -4700
rect 3830 -4710 4030 -4690
rect 3830 -4880 3850 -4710
rect 4010 -4840 4030 -4710
rect 4101 -4719 4300 -4686
rect 3831 -5160 3850 -4880
rect 3830 -5330 3850 -5160
rect 3830 -5350 3851 -5330
rect 3360 -5850 3760 -5830
rect 3831 -5830 3851 -5350
rect 4011 -5830 4030 -4840
rect 3831 -5850 4030 -5830
rect 4100 -4720 4300 -4719
rect 4100 -5830 4120 -4720
rect 4280 -4725 4300 -4720
rect 4370 -4710 4570 -4690
rect 4280 -5360 4299 -4725
rect 4370 -4880 4390 -4710
rect 4550 -4781 4570 -4710
rect 4371 -5160 4390 -4880
rect 4370 -5330 4390 -5160
rect 4551 -4880 4570 -4781
rect 4551 -5160 4569 -4880
rect 4370 -5350 4391 -5330
rect 4280 -5830 4300 -5360
rect 4100 -5850 4300 -5830
rect 4371 -5831 4391 -5350
rect 4551 -5831 4570 -5160
rect 4371 -5851 4570 -5831
rect 220 -6030 830 -6020
rect 220 -6130 240 -6030
rect 810 -6130 830 -6030
rect 220 -6150 830 -6130
rect -990 -6200 -380 -6180
rect -990 -6300 -970 -6200
rect -400 -6300 -380 -6200
rect -990 -6320 -380 -6300
<< viali >>
rect -3780 -1210 4640 -900
rect -970 -2000 -400 -1900
rect 240 -2000 810 -1900
rect -3780 -2760 -3630 -2221
rect -3580 -2760 -3430 -2221
rect -3290 -2750 -2770 -2230
rect -3290 -2970 -2770 -2900
rect -3780 -4230 -3630 -3100
rect -3580 -4230 -3430 -3100
rect -3309 -4233 -3157 -3106
rect -3041 -4230 -3040 -3111
rect -3040 -4230 -2890 -3111
rect -2890 -4230 -2889 -3111
rect -3041 -4234 -2889 -4230
rect -2770 -4232 -2618 -3105
rect -2504 -3110 -2352 -3109
rect -2504 -4230 -2500 -3110
rect -2500 -4230 -2352 -3110
rect -2504 -4232 -2352 -4230
rect -2234 -4228 -2230 -3101
rect -2230 -4228 -2082 -3101
rect -1360 -3250 -1230 -2120
rect -1140 -3250 -1010 -2120
rect -880 -3250 -750 -2120
rect -610 -3250 -480 -2120
rect -360 -3250 -230 -2120
rect -130 -3240 -30 -2140
rect 60 -3250 190 -2120
rect 320 -3250 450 -2120
rect 590 -3240 720 -2110
rect 850 -3240 980 -2110
rect 1080 -3250 1210 -2120
rect 2690 -2130 4340 -2040
rect 2290 -2410 2440 -2250
rect 2490 -2410 2650 -2250
rect 1360 -3290 1450 -3200
rect 2300 -3220 2427 -2410
rect 2290 -3380 2440 -3220
rect 2497 -3355 2635 -2410
rect 2758 -3063 2916 -2279
rect 2759 -3384 2915 -3063
rect 3037 -3027 3195 -2277
rect 3036 -3063 3195 -3027
rect 3036 -3379 3192 -3063
rect 3300 -3063 3458 -2281
rect 3301 -3393 3457 -3063
rect 3569 -3045 3727 -2287
rect 3569 -3063 3728 -3045
rect 3572 -3397 3728 -3063
rect 3841 -3038 3999 -2282
rect 3838 -3063 3999 -3038
rect 3838 -3390 3994 -3063
rect 4114 -3045 4272 -2277
rect 4114 -3063 4274 -3045
rect 4118 -3397 4274 -3063
rect 4382 -3031 4540 -2279
rect 4680 -2410 4832 -2250
rect 4381 -3063 4540 -3031
rect 4381 -3383 4537 -3063
rect 4682 -3369 4832 -2410
rect -430 -3640 -40 -3560
rect -900 -4250 -740 -3730
rect -700 -4250 -540 -3730
rect 1360 -3690 1450 -3600
rect -430 -4250 -270 -3730
rect -160 -4250 0 -3730
rect 110 -4250 270 -3730
rect 380 -4250 540 -3730
rect 590 -4250 750 -3730
rect -3290 -4990 -1780 -4400
rect 380 -4520 730 -4390
rect 2370 -4440 2960 -4020
rect 4370 -4260 4730 -3900
rect 2370 -4480 3670 -4440
rect 2370 -4560 3400 -4480
rect 2370 -4600 2720 -4560
rect 2720 -4590 3400 -4560
rect 3400 -4590 3670 -4480
rect 2720 -4600 3670 -4590
rect -1360 -5920 -1230 -4790
rect -1140 -5920 -1010 -4790
rect -880 -5920 -750 -4790
rect -610 -5920 -480 -4790
rect -360 -5920 -230 -4790
rect -130 -5910 -30 -4810
rect 60 -5920 190 -4790
rect 320 -5920 450 -4790
rect 590 -5910 720 -4780
rect 850 -5910 980 -4780
rect 1080 -5920 1210 -4790
rect 2930 -5400 2990 -5150
rect 2350 -5940 2690 -5510
rect 3380 -5830 3540 -4700
rect 3580 -5830 3740 -4700
rect 3850 -4840 4010 -4710
rect 3850 -5330 4011 -4840
rect 3851 -5830 4011 -5330
rect 4120 -5830 4280 -4720
rect 4390 -4781 4550 -4710
rect 4390 -5330 4551 -4781
rect 4391 -5831 4551 -5330
rect 240 -6130 810 -6030
rect -970 -6300 -400 -6200
rect -3770 -6800 4650 -6470
rect -3120 -7360 4170 -7060
<< metal1 >>
rect -3900 -900 4680 -860
rect -3900 -1210 -3780 -900
rect 4640 -1210 4680 -900
rect -3900 -1250 4680 -1210
rect -3900 -1820 4330 -1370
rect -3810 -2221 -3420 -2190
rect -3810 -2760 -3780 -2221
rect -3630 -2760 -3580 -2221
rect -3430 -2760 -3420 -2221
rect -3810 -3050 -3420 -2760
rect -3330 -2230 -2730 -1820
rect -3330 -2750 -3290 -2230
rect -2770 -2750 -2730 -2230
rect -3330 -2900 -2730 -2750
rect -3330 -2970 -3290 -2900
rect -2770 -2970 -2730 -2900
rect -3330 -3010 -2730 -2970
rect -1590 -1900 -380 -1880
rect -1590 -2000 -970 -1900
rect -400 -2000 -380 -1900
rect -1590 -2020 -380 -2000
rect 220 -1900 1470 -1880
rect 220 -2000 240 -1900
rect 810 -2000 1470 -1900
rect 220 -2020 1470 -2000
rect -3820 -3100 -3420 -3050
rect -3820 -3290 -3780 -3100
rect -3810 -4230 -3780 -3290
rect -3630 -4230 -3580 -3100
rect -3430 -3690 -3420 -3100
rect -3329 -3106 -3130 -3088
rect -3430 -3920 -3402 -3690
rect -3430 -4230 -3420 -3920
rect -3329 -4201 -3309 -3106
rect -3810 -4260 -3420 -4230
rect -3330 -4233 -3309 -4201
rect -3157 -4233 -3130 -3106
rect -3330 -4253 -3130 -4233
rect -3059 -3111 -2859 -3091
rect -3059 -4234 -3041 -3111
rect -2889 -4234 -2859 -3111
rect -2790 -3105 -2591 -3087
rect -2790 -4177 -2770 -3105
rect -3330 -4330 -3131 -4253
rect -3059 -4254 -2859 -4234
rect -2791 -4232 -2770 -4177
rect -2618 -4232 -2591 -3105
rect -2791 -4252 -2591 -4232
rect -2518 -3109 -2318 -3091
rect -2518 -4232 -2504 -3109
rect -2352 -4232 -2318 -3109
rect -2248 -3101 -2050 -3091
rect -2248 -4155 -2234 -3101
rect -2791 -4330 -2592 -4252
rect -2518 -4254 -2318 -4232
rect -2249 -4228 -2234 -4155
rect -2082 -4228 -2050 -3101
rect -2249 -4330 -2050 -4228
rect -1985 -4266 -1777 -3084
rect -1953 -4330 -1710 -4329
rect -3360 -4400 -1710 -4330
rect -3360 -4990 -3290 -4400
rect -1780 -4990 -1710 -4400
rect -3360 -5040 -1710 -4990
rect -1590 -5920 -1460 -2020
rect -1390 -2120 -1210 -2090
rect -1390 -3250 -1360 -2120
rect -1230 -3250 -1210 -2120
rect -1390 -3270 -1210 -3250
rect -1170 -2120 -990 -2090
rect -1170 -3250 -1140 -2120
rect -1010 -3250 -990 -2120
rect -1170 -3270 -990 -3250
rect -910 -2120 -730 -2090
rect -910 -3250 -880 -2120
rect -750 -3250 -730 -2120
rect -910 -3340 -730 -3250
rect -640 -2120 -460 -2090
rect -640 -3250 -610 -2120
rect -480 -3250 -460 -2120
rect -640 -3270 -460 -3250
rect -380 -2120 -200 -2090
rect -380 -3250 -360 -2120
rect -230 -3250 -200 -2120
rect -380 -3340 -200 -3250
rect -150 -2140 -10 -2110
rect -150 -3240 -130 -2140
rect -30 -3240 -10 -2140
rect -150 -3260 -10 -3240
rect 40 -2120 220 -2090
rect 40 -3250 60 -2120
rect 190 -3250 220 -2120
rect -910 -3530 -200 -3340
rect 40 -3360 220 -3250
rect 300 -2120 480 -2090
rect 300 -3250 320 -2120
rect 450 -3250 480 -2120
rect 570 -2110 750 -2090
rect 570 -3030 590 -2110
rect 300 -3270 480 -3250
rect 560 -3240 590 -3030
rect 720 -3240 750 -2110
rect 560 -3270 750 -3240
rect 830 -2110 1010 -2090
rect 830 -3240 850 -2110
rect 980 -3240 1010 -2110
rect 830 -3270 1010 -3240
rect 1050 -2120 1230 -2090
rect 1050 -3250 1080 -2120
rect 1210 -3250 1230 -2120
rect 1050 -3270 1230 -3250
rect 1340 -3200 1470 -2020
rect 2670 -1990 4330 -1820
rect 2670 -2040 4360 -1990
rect 2670 -2130 2690 -2040
rect 4340 -2130 4360 -2040
rect 2670 -2150 4360 -2130
rect 2273 -2230 2654 -2228
rect 2270 -2250 2669 -2230
rect 2270 -2410 2290 -2250
rect 2440 -2410 2490 -2250
rect 2650 -2410 2669 -2250
rect 2270 -2430 2300 -2410
rect 2273 -3200 2300 -2430
rect 560 -3360 740 -3270
rect 1340 -3290 1360 -3200
rect 1450 -3290 1470 -3200
rect 1340 -3300 1470 -3290
rect 2270 -3220 2300 -3200
rect 2427 -3220 2497 -2410
rect 40 -3510 2020 -3360
rect 2270 -3380 2290 -3220
rect 2440 -3355 2497 -3220
rect 2635 -2430 2669 -2410
rect 2745 -2279 2933 -2224
rect 2635 -3355 2654 -2430
rect 2745 -3016 2758 -2279
rect 2440 -3380 2654 -3355
rect 2270 -3400 2654 -3380
rect 2741 -3063 2758 -3016
rect 2916 -3016 2933 -2279
rect 3016 -2277 3204 -2227
rect 3016 -2280 3037 -2277
rect 3195 -2280 3204 -2277
rect 3016 -3016 3030 -2280
rect 2916 -3063 2938 -3016
rect 2741 -3384 2759 -3063
rect 2915 -3262 2938 -3063
rect 2915 -3384 2939 -3262
rect -90 -3530 -8 -3529
rect -910 -3560 -8 -3530
rect -910 -3620 -430 -3560
rect -450 -3640 -430 -3620
rect -40 -3640 -8 -3560
rect -450 -3647 -8 -3640
rect 100 -3550 2020 -3510
rect 2741 -3515 2939 -3384
rect 3013 -3380 3030 -3016
rect 3200 -3016 3204 -2280
rect 3286 -2281 3474 -2222
rect 3200 -3380 3210 -3016
rect 3286 -3020 3300 -2281
rect 3282 -3063 3300 -3020
rect 3458 -3020 3474 -2281
rect 3555 -2287 3743 -2233
rect 3555 -3015 3569 -2287
rect 3458 -3063 3479 -3020
rect 3282 -3369 3301 -3063
rect 3013 -3409 3210 -3380
rect 3281 -3393 3301 -3369
rect 3457 -3393 3479 -3063
rect 3281 -3515 3479 -3393
rect 3550 -3063 3569 -3015
rect 3550 -3397 3572 -3063
rect 3727 -3015 3743 -2287
rect 3826 -2282 4014 -2233
rect 3826 -3015 3841 -2282
rect 3727 -3045 3747 -3015
rect 3728 -3397 3747 -3045
rect 3550 -3408 3747 -3397
rect 3820 -3038 3841 -3015
rect 3999 -3015 4014 -2282
rect 4100 -2277 4288 -2234
rect 3820 -3390 3838 -3038
rect 3999 -3063 4017 -3015
rect 4100 -3017 4114 -2277
rect 3994 -3358 4017 -3063
rect 4092 -3063 4114 -3017
rect 3994 -3390 4018 -3358
rect 3820 -3515 4018 -3390
rect 4092 -3397 4118 -3063
rect 4272 -3017 4288 -2277
rect 4363 -2279 4551 -2233
rect 4272 -3045 4289 -3017
rect 4274 -3397 4289 -3045
rect 4363 -3031 4382 -2279
rect 4540 -3015 4551 -2279
rect 4660 -2250 4860 -2230
rect 4660 -2410 4680 -2250
rect 4660 -2430 4682 -2410
rect 4363 -3301 4381 -3031
rect 4540 -3063 4560 -3015
rect 4092 -3410 4289 -3397
rect 4362 -3383 4381 -3301
rect 4537 -3383 4560 -3063
rect 4362 -3515 4560 -3383
rect 4663 -3369 4682 -2430
rect 4832 -3369 4860 -2250
rect 4663 -3406 4860 -3369
rect 2709 -3520 4567 -3515
rect 100 -3600 1240 -3550
rect 1340 -3600 1470 -3590
rect -450 -3650 -10 -3647
rect -920 -3730 -530 -3710
rect -920 -4250 -900 -3730
rect -740 -4250 -700 -3730
rect -540 -4250 -530 -3730
rect -450 -3730 -250 -3650
rect -450 -3770 -430 -3730
rect -441 -3905 -430 -3770
rect -920 -4270 -530 -4250
rect -440 -4250 -430 -3905
rect -270 -3770 -250 -3730
rect -170 -3730 10 -3710
rect -270 -3905 -254 -3770
rect -270 -4250 -260 -3905
rect -440 -4270 -260 -4250
rect -170 -4250 -160 -3730
rect 0 -4250 10 -3730
rect -170 -4270 10 -4250
rect 100 -3730 280 -3600
rect 1340 -3690 1360 -3600
rect 1450 -3690 1470 -3600
rect 100 -4250 110 -3730
rect 270 -4250 280 -3730
rect 100 -4310 280 -4250
rect 370 -3730 760 -3710
rect 370 -4250 380 -3730
rect 540 -4250 590 -3730
rect 750 -4250 760 -3730
rect 370 -4270 760 -4250
rect -910 -4490 280 -4310
rect 340 -4390 770 -4350
rect -910 -4640 -200 -4490
rect 340 -4520 380 -4390
rect 730 -4520 770 -4390
rect 340 -4540 770 -4520
rect -3900 -6020 -1460 -5920
rect -1390 -4790 -1210 -4760
rect -1390 -5920 -1360 -4790
rect -1230 -5920 -1210 -4790
rect -1390 -5940 -1210 -5920
rect -1170 -4790 -990 -4760
rect -1170 -5920 -1140 -4790
rect -1010 -5920 -990 -4790
rect -1170 -5940 -990 -5920
rect -910 -4790 -730 -4640
rect -910 -5920 -880 -4790
rect -750 -5920 -730 -4790
rect -910 -5950 -730 -5920
rect -640 -4790 -460 -4760
rect -640 -5920 -610 -4790
rect -480 -5920 -460 -4790
rect -640 -5940 -460 -5920
rect -380 -4790 -200 -4640
rect 40 -4680 770 -4540
rect -380 -5920 -360 -4790
rect -230 -5920 -200 -4790
rect -380 -5950 -200 -5920
rect -150 -4810 -10 -4780
rect -150 -5910 -130 -4810
rect -30 -5910 -10 -4810
rect -150 -5930 -10 -5910
rect 40 -4790 220 -4680
rect 40 -5920 60 -4790
rect 190 -5920 220 -4790
rect 40 -5950 220 -5920
rect 300 -4790 480 -4760
rect 300 -5920 320 -4790
rect 450 -5920 480 -4790
rect 570 -4780 750 -4680
rect 570 -5700 590 -4780
rect 300 -5940 480 -5920
rect 560 -5910 590 -5700
rect 720 -5910 750 -4780
rect 560 -5940 750 -5910
rect 830 -4780 1010 -4760
rect 830 -5910 850 -4780
rect 980 -5910 1010 -4780
rect 830 -5940 1010 -5910
rect 1050 -4790 1230 -4760
rect 1050 -5920 1080 -4790
rect 1210 -5920 1230 -4790
rect 1050 -5940 1230 -5920
rect 560 -5950 740 -5940
rect -3900 -6030 830 -6020
rect -3900 -6060 240 -6030
rect -1590 -6130 240 -6060
rect 810 -6130 830 -6030
rect -1590 -6150 830 -6130
rect 1340 -6180 1470 -3690
rect 1590 -3980 2020 -3550
rect 2450 -3625 4567 -3520
rect 2450 -3880 4570 -3625
rect 2450 -3898 4830 -3880
rect 2450 -3900 2850 -3898
rect 3133 -3900 4830 -3898
rect 1590 -4020 2990 -3980
rect 1590 -4440 2370 -4020
rect 2960 -4420 2990 -4020
rect 3133 -4260 4370 -3900
rect 4730 -4260 4830 -3900
rect 3133 -4280 4830 -4260
rect 3133 -4285 4570 -4280
rect 3133 -4287 3736 -4285
rect 3133 -4290 3629 -4287
rect 3830 -4360 4570 -4285
rect 2960 -4440 3730 -4420
rect 2320 -4600 2370 -4440
rect 3670 -4600 3730 -4440
rect 2320 -4610 3730 -4600
rect 3350 -4679 3560 -4670
rect 3350 -4680 3603 -4679
rect 3350 -4700 3760 -4680
rect 2900 -5150 3020 -5120
rect 2900 -5400 2930 -5150
rect 2990 -5400 3020 -5150
rect 2900 -5430 3020 -5400
rect 2320 -5510 2720 -5470
rect 2320 -5940 2350 -5510
rect 2690 -5940 2720 -5510
rect 2320 -5980 2720 -5940
rect -3890 -6200 1470 -6180
rect -3890 -6300 -970 -6200
rect -400 -6300 1470 -6200
rect -3890 -6310 1470 -6300
rect -3890 -6320 1350 -6310
rect 2910 -6430 3010 -5430
rect 3350 -5830 3380 -4700
rect 3540 -5830 3580 -4700
rect 3740 -5830 3760 -4700
rect 3830 -4710 4030 -4360
rect 3830 -5330 3850 -4710
rect 4010 -4840 4030 -4710
rect 4101 -4719 4300 -4686
rect 3830 -5350 3851 -5330
rect 3350 -6430 3760 -5830
rect 3831 -5830 3851 -5350
rect 4011 -5830 4030 -4840
rect 3831 -5850 4030 -5830
rect 4100 -4720 4300 -4719
rect 4100 -5830 4120 -4720
rect 4280 -4725 4300 -4720
rect 4370 -4710 4570 -4360
rect 4280 -5370 4299 -4725
rect 4370 -5330 4390 -4710
rect 4550 -4781 4570 -4710
rect 4370 -5350 4391 -5330
rect 4280 -5830 4300 -5370
rect 4100 -6430 4300 -5830
rect 4371 -5831 4391 -5350
rect 4551 -5831 4570 -4781
rect 4371 -5851 4570 -5831
rect -3910 -6470 4690 -6430
rect -3910 -6800 -3770 -6470
rect 4650 -6800 4690 -6470
rect -3910 -6840 4690 -6800
rect -3230 -7060 4270 -6840
rect -3230 -7360 -3120 -7060
rect 4170 -7360 4270 -7060
rect -3230 -7450 4270 -7360
<< via1 >>
rect -3780 -1210 4640 -900
rect -3780 -2760 -3630 -2221
rect -3580 -2760 -3430 -2221
rect -3780 -4230 -3630 -3100
rect -3580 -4230 -3430 -3100
rect -3041 -4234 -2889 -3111
rect -2504 -4232 -2352 -3109
rect -3290 -4990 -1780 -4400
rect -1360 -3250 -1230 -2120
rect -1140 -3250 -1010 -2120
rect -610 -3250 -480 -2120
rect -130 -3240 -30 -2140
rect 320 -3250 450 -2120
rect 850 -3240 980 -2110
rect 1080 -3250 1210 -2120
rect 2290 -2410 2440 -2250
rect 2490 -2410 2650 -2250
rect 1360 -3290 1450 -3200
rect 2300 -3220 2427 -2410
rect 2290 -3380 2440 -3220
rect 2497 -3355 2635 -2410
rect 3030 -3027 3037 -2280
rect 3037 -3027 3195 -2280
rect 3030 -3379 3036 -3027
rect 3036 -3063 3195 -3027
rect 3195 -3063 3200 -2280
rect 3036 -3379 3192 -3063
rect 3192 -3379 3200 -3063
rect 3030 -3380 3200 -3379
rect 3580 -3390 3720 -2290
rect 4120 -3390 4260 -2290
rect 4680 -2410 4832 -2250
rect 4682 -3369 4832 -2410
rect -900 -4250 -740 -3730
rect -700 -4250 -540 -3730
rect -160 -4250 0 -3730
rect 1360 -3690 1450 -3600
rect 380 -4250 540 -3730
rect 590 -4250 750 -3730
rect -1360 -5920 -1230 -4790
rect -1140 -5920 -1010 -4790
rect -610 -5920 -480 -4790
rect -130 -5910 -30 -4810
rect 320 -5920 450 -4790
rect 850 -5910 980 -4780
rect 1080 -5920 1210 -4790
rect 4370 -4260 4730 -3900
rect 2350 -5940 2690 -5510
rect -3770 -6800 4650 -6470
rect -3120 -7360 4170 -7060
<< metal2 >>
rect -3810 -900 4860 -860
rect -3810 -1210 -3780 -900
rect 4640 -1210 4860 -900
rect -3810 -1250 4860 -1210
rect -3810 -2221 -3410 -1250
rect -3810 -2760 -3780 -2221
rect -3630 -2760 -3580 -2221
rect -3430 -2760 -3410 -2221
rect -3810 -3068 -3410 -2760
rect -1390 -2120 -1210 -2090
rect -3810 -3100 -1750 -3068
rect -3810 -4230 -3780 -3100
rect -3630 -4230 -3580 -3100
rect -3430 -3109 -1750 -3100
rect -3430 -3111 -2504 -3109
rect -3430 -4230 -3041 -3111
rect -3810 -4234 -3041 -4230
rect -2889 -4232 -2504 -3111
rect -2352 -4232 -1750 -3109
rect -1390 -3250 -1360 -2120
rect -1230 -3250 -1210 -2120
rect -1170 -2120 -990 -2090
rect -1170 -3160 -1140 -2120
rect -1390 -3270 -1210 -3250
rect -1180 -3250 -1140 -3160
rect -1010 -3250 -990 -2120
rect -1180 -3360 -990 -3250
rect -640 -2120 -460 -2090
rect -640 -3250 -610 -2120
rect -480 -3250 -460 -2120
rect -640 -3360 -460 -3250
rect -150 -2140 -10 -2110
rect -150 -3240 -130 -2140
rect -30 -3240 -10 -2140
rect -150 -3260 -10 -3240
rect 300 -2120 480 -2090
rect 300 -3250 320 -2120
rect 450 -3250 480 -2120
rect 300 -3360 480 -3250
rect 830 -2110 1010 -2090
rect 830 -3240 850 -2110
rect 980 -3240 1010 -2110
rect 830 -3360 1010 -3240
rect 1050 -2120 1230 -2090
rect 1050 -3250 1080 -2120
rect 1210 -3250 1230 -2120
rect 2270 -2250 4860 -1250
rect 2270 -2410 2290 -2250
rect 2440 -2410 2490 -2250
rect 2650 -2280 4680 -2250
rect 2650 -2410 3030 -2280
rect 1050 -3270 1230 -3250
rect 1350 -3200 1460 -3190
rect -1410 -3370 1010 -3360
rect -2889 -4234 -1750 -4232
rect -3810 -4264 -1750 -4234
rect -1630 -3650 1010 -3370
rect 1350 -3290 1360 -3200
rect 1450 -3290 1460 -3200
rect 1350 -3600 1460 -3290
rect 2270 -3220 2300 -2410
rect 2427 -3220 2497 -2410
rect 2270 -3380 2290 -3220
rect 2440 -3355 2497 -3220
rect 2635 -3355 3030 -2410
rect 2440 -3380 3030 -3355
rect 3200 -2290 4680 -2280
rect 3200 -3380 3580 -2290
rect 2270 -3390 3580 -3380
rect 3720 -3390 4120 -2290
rect 4260 -2410 4680 -2290
rect 4260 -3369 4682 -2410
rect 4832 -3369 4860 -2250
rect 4260 -3390 4860 -3369
rect 2270 -3400 4860 -3390
rect 2270 -3401 2667 -3400
rect 3011 -3416 3208 -3400
rect 3556 -3408 3753 -3400
rect 4093 -3413 4290 -3400
rect 4663 -3406 4860 -3400
rect -3810 -4280 -3410 -4264
rect -1985 -4266 -1777 -4264
rect -1630 -4330 -1380 -3650
rect 1350 -3690 1360 -3600
rect 1450 -3690 1460 -3600
rect 1350 -3700 1460 -3690
rect -920 -3730 -530 -3710
rect -920 -3740 -900 -3730
rect -1010 -4240 -900 -3740
rect -920 -4250 -900 -4240
rect -740 -4250 -700 -3730
rect -540 -3740 -530 -3730
rect -170 -3730 10 -3710
rect -170 -3740 -160 -3730
rect -540 -4240 -160 -3740
rect -540 -4250 -530 -4240
rect -920 -4270 -530 -4250
rect -170 -4250 -160 -4240
rect 0 -3740 10 -3730
rect 370 -3730 760 -3710
rect 370 -3740 380 -3730
rect 0 -4240 380 -3740
rect 0 -4250 10 -4240
rect -170 -4270 10 -4250
rect 370 -4250 380 -4240
rect 540 -4250 590 -3730
rect 750 -3740 760 -3730
rect 750 -4240 1650 -3740
rect 750 -4250 760 -4240
rect 370 -4270 760 -4250
rect -3360 -4400 1030 -4330
rect -3360 -4990 -3290 -4400
rect -1780 -4620 1030 -4400
rect -1780 -4660 1010 -4620
rect -1780 -4990 -1450 -4660
rect -3360 -5040 -1450 -4990
rect -1390 -4790 -1210 -4760
rect -1390 -5920 -1360 -4790
rect -1230 -5920 -1210 -4790
rect -1170 -4790 -990 -4660
rect -1170 -5830 -1140 -4790
rect -1390 -5940 -1210 -5920
rect -1180 -5920 -1140 -5830
rect -1010 -5920 -990 -4790
rect -1180 -5950 -990 -5920
rect -640 -4790 -460 -4660
rect -640 -5920 -610 -4790
rect -480 -5920 -460 -4790
rect -640 -5950 -460 -5920
rect -150 -4810 -10 -4780
rect -150 -5910 -130 -4810
rect -30 -5910 -10 -4810
rect -150 -5930 -10 -5910
rect 300 -4790 480 -4660
rect 300 -5920 320 -4790
rect 450 -5920 480 -4790
rect 300 -5950 480 -5920
rect 830 -4780 1010 -4660
rect 830 -5910 850 -4780
rect 980 -5910 1010 -4780
rect 830 -5950 1010 -5910
rect 1050 -4790 1230 -4760
rect 1050 -5920 1080 -4790
rect 1210 -5920 1230 -4790
rect 1050 -5940 1230 -5920
rect 1330 -6430 1650 -4240
rect 4350 -3900 4750 -3880
rect 4350 -4260 4370 -3900
rect 4730 -4260 4750 -3900
rect 4350 -4280 4750 -4260
rect 2320 -5510 2720 -5470
rect 2320 -5940 2350 -5510
rect 2690 -5940 2720 -5510
rect 2320 -5980 2720 -5940
rect -3800 -6470 4690 -6430
rect -3800 -6800 -3770 -6470
rect 4650 -6800 4690 -6470
rect -3800 -6840 4690 -6800
rect -3230 -7060 4270 -6840
rect -3230 -7360 -3120 -7060
rect 4170 -7360 4270 -7060
rect -3230 -7450 4270 -7360
<< via2 >>
rect -3780 -1210 4640 -900
rect -1360 -3250 -1230 -2120
rect -130 -3240 -30 -2140
rect 1080 -3250 1210 -2120
rect -1360 -5920 -1230 -4790
rect -130 -5910 -30 -4810
rect 1080 -5920 1210 -4790
rect 4370 -4260 4730 -3900
rect 2350 -5940 2690 -5510
rect -3770 -6800 4650 -6470
rect -3120 -7360 4170 -7060
<< metal3 >>
rect -3810 -900 4680 -860
rect -3810 -1210 -3780 -900
rect 4640 -1210 4680 -900
rect -3810 -1250 4680 -1210
rect -1670 -2120 -1180 -1250
rect -1670 -3250 -1360 -2120
rect -1230 -3250 -1180 -2120
rect -1670 -4790 -1180 -3250
rect -1670 -5920 -1360 -4790
rect -1230 -5920 -1180 -4790
rect -1670 -6080 -1180 -5920
rect -320 -2140 170 -1250
rect -320 -3240 -130 -2140
rect -30 -3240 170 -2140
rect -320 -4810 170 -3240
rect -320 -5910 -130 -4810
rect -30 -5910 170 -4810
rect -320 -6100 170 -5910
rect 1030 -2120 1530 -1250
rect 1030 -3250 1080 -2120
rect 1210 -3250 1530 -2120
rect 1030 -4790 1530 -3250
rect 1030 -5920 1080 -4790
rect 1210 -5920 1530 -4790
rect 2030 -3880 4120 -3030
rect 2030 -3900 4750 -3880
rect 2030 -4260 4370 -3900
rect 4730 -4260 4750 -3900
rect 2030 -4290 4750 -4260
rect 2030 -5120 4120 -4290
rect 1030 -6050 1530 -5920
rect 2320 -5510 2720 -5470
rect 2320 -5940 2350 -5510
rect 2690 -5940 2720 -5510
rect 2320 -5980 2720 -5940
rect 1040 -6090 1530 -6050
rect -3800 -6470 4690 -6430
rect -3800 -6800 -3770 -6470
rect 4650 -6800 4690 -6470
rect -3800 -6840 4690 -6800
rect -3230 -7060 4270 -6840
rect -3230 -7360 -3120 -7060
rect 4170 -7360 4270 -7060
rect -3230 -7450 4270 -7360
<< via3 >>
rect 2350 -5940 2690 -5510
<< mimcap >>
rect 2070 -3790 4070 -3080
rect 2070 -4290 2320 -3790
rect 2820 -4290 4070 -3790
rect 2070 -5080 4070 -4290
<< mimcapcontact >>
rect 2320 -4290 2820 -3790
<< metal4 >>
rect -5040 -750 5960 250
rect -5040 -6950 -4040 -750
rect 2280 -3790 2860 -3720
rect 2280 -4290 2320 -3790
rect 2820 -4290 2860 -3790
rect 2280 -5510 2860 -4290
rect 4960 -5160 5960 -750
rect 2280 -5940 2350 -5510
rect 2690 -5940 2860 -5510
rect 2280 -6010 2860 -5940
rect 5030 -6220 5960 -5160
rect 5010 -6230 5960 -6220
rect -3230 -6950 4270 -6540
rect 4960 -6950 5960 -6230
rect -5040 -7060 5960 -6950
rect -5040 -7360 -3120 -7060
rect 4170 -7360 5960 -7060
rect -5040 -7950 5960 -7360
<< via4 >>
rect -3120 -7360 4170 -7060
<< metal5 >>
rect -5040 -750 5960 250
rect -5040 -6950 -4040 -750
rect -3230 -6950 4270 -6540
rect 4960 -6950 5960 -750
rect -5040 -7060 5960 -6950
rect -5040 -7360 -3120 -7060
rect 4170 -7360 5960 -7060
rect -5040 -7950 5960 -7360
<< labels >>
rlabel metal1 -3900 -1160 -3900 -1160 7 VDD
port 1 w
rlabel metal1 -3900 -1650 -3900 -1650 7 Bias1
port 3 w
rlabel metal1 4830 -4080 4830 -4080 3 OUT
port 2 e
rlabel metal1 -3900 -5990 -3900 -5990 7 INN
port 5 w
rlabel metal1 -3890 -6260 -3890 -6260 1 INP
port 4 n
rlabel metal1 -3910 -6750 -3910 -6750 7 VSS
port 6 w
<< end >>
